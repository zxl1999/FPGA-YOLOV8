// megafunction wizard: %FIFO%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: dcfifo_mixed_widths 

// ============================================================
// File Name: cmos1_fifo.v
// Megafunction Name(s):
// 			dcfifo_mixed_widths
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.1.0 Build 162 10/23/2013 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module cmos1_fifo (
	aclr,
	data,
	rdclk,
	rdreq,
	wrclk,
	wrreq,
	q,
	rdempty,
	rdusedw,
	wrfull,
	wrusedw);

	input	  aclr;
	input	[7:0]  data;
	input	  rdclk;
	input	  rdreq;
	input	  wrclk;
	input	  wrreq;
	output reg [31:0]  q;
	output	  rdempty;
	output	[9:0]  rdusedw;
	output	  wrfull;
	output	[11:0]  wrusedw;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri0	  aclr;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [31:0] sub_wire1;
	wire  sub_wire2;
	wire [11:0] sub_wire3;
	wire [9:0] sub_wire4;
	wire  wrfull = sub_wire0;
	
	wire  rdempty = sub_wire2;
	wire [11:0] wrusedw = sub_wire3[11:0];
	wire [9:0] rdusedw = sub_wire4[9:0];
	
	always @(posedge rdclk) begin
	q = sub_wire1[31:0];
    if (rdreq && !rdempty) begin
		q[0] = (sub_wire1[31] & 1'b1) ^ (sub_wire1[0] & 1'b1) ^ (sub_wire1[1] & 1'b1);
q[1] = (sub_wire1[0] & 1'b1) ^ (sub_wire1[1] & 1'b1) ^ (sub_wire1[2] & 1'b1);
q[2] = (sub_wire1[1] & 1'b1) ^ (sub_wire1[2] & 1'b1) ^ (sub_wire1[3] & 1'b1);
q[3] = (sub_wire1[2] & 1'b1) ^ (sub_wire1[3] & 1'b1) ^ (sub_wire1[4] & 1'b1);
q[4] = (sub_wire1[3] & 1'b1) ^ (sub_wire1[4] & 1'b1) ^ (sub_wire1[5] & 1'b1);
q[5] = (sub_wire1[4] & 1'b1) ^ (sub_wire1[5] & 1'b1) ^ (sub_wire1[6] & 1'b1);
q[6] = (sub_wire1[5] & 1'b1) ^ (sub_wire1[6] & 1'b1) ^ (sub_wire1[7] & 1'b1);
q[7] = (sub_wire1[6] & 1'b1) ^ (sub_wire1[7] & 1'b1) ^ (sub_wire1[8] & 1'b1);
q[8] = (sub_wire1[7] & 1'b1) ^ (sub_wire1[8] & 1'b1) ^ (sub_wire1[9] & 1'b1);
q[9] = (sub_wire1[8] & 1'b1) ^ (sub_wire1[9] & 1'b1) ^ (sub_wire1[10] & 1'b1);
q[10] = (sub_wire1[9] & 1'b1) ^ (sub_wire1[10] & 1'b1) ^ (sub_wire1[11] & 1'b1);
q[11] = (sub_wire1[10] & 1'b1) ^ (sub_wire1[11] & 1'b1) ^ (sub_wire1[12] & 1'b1);
q[12] = (sub_wire1[11] & 1'b1) ^ (sub_wire1[12] & 1'b1) ^ (sub_wire1[13] & 1'b1);
q[13] = (sub_wire1[12] & 1'b1) ^ (sub_wire1[13] & 1'b1) ^ (sub_wire1[14] & 1'b1);
q[14] = (sub_wire1[13] & 1'b1) ^ (sub_wire1[14] & 1'b1) ^ (sub_wire1[15] & 1'b1);
q[15] = (sub_wire1[14] & 1'b1) ^ (sub_wire1[15] & 1'b1) ^ (sub_wire1[16] & 1'b1);
q[16] = (sub_wire1[15] & 1'b1) ^ (sub_wire1[16] & 1'b1) ^ (sub_wire1[17] & 1'b1);
q[17] = (sub_wire1[16] & 1'b1) ^ (sub_wire1[17] & 1'b1) ^ (sub_wire1[18] & 1'b1);
q[18] = (sub_wire1[17] & 1'b1) ^ (sub_wire1[18] & 1'b1) ^ (sub_wire1[19] & 1'b1);
q[19] = (sub_wire1[18] & 1'b1) ^ (sub_wire1[19] & 1'b1) ^ (sub_wire1[20] & 1'b1);
q[20] = (sub_wire1[19] & 1'b1) ^ (sub_wire1[20] & 1'b1) ^ (sub_wire1[21] & 1'b1);
q[21] = (sub_wire1[20] & 1'b1) ^ (sub_wire1[21] & 1'b1) ^ (sub_wire1[22] & 1'b1);
q[22] = (sub_wire1[21] & 1'b1) ^ (sub_wire1[22] & 1'b1) ^ (sub_wire1[23] & 1'b1);
q[23] = (sub_wire1[22] & 1'b1) ^ (sub_wire1[23] & 1'b1) ^ (sub_wire1[24] & 1'b1);
q[24] = (sub_wire1[23] & 1'b1) ^ (sub_wire1[24] & 1'b1) ^ (sub_wire1[25] & 1'b1);
q[25] = (sub_wire1[24] & 1'b1) ^ (sub_wire1[25] & 1'b1) ^ (sub_wire1[26] & 1'b1);
q[26] = (sub_wire1[25] & 1'b1) ^ (sub_wire1[26] & 1'b1) ^ (sub_wire1[27] & 1'b1);
q[27] = (sub_wire1[26] & 1'b1) ^ (sub_wire1[27] & 1'b1) ^ (sub_wire1[28] & 1'b1);
q[28] = (sub_wire1[27] & 1'b1) ^ (sub_wire1[28] & 1'b1) ^ (sub_wire1[29] & 1'b1);
q[29] = (sub_wire1[28] & 1'b1) ^ (sub_wire1[29] & 1'b1) ^ (sub_wire1[30] & 1'b1);
q[30] = (sub_wire1[29] & 1'b1) ^ (sub_wire1[30] & 1'b1) ^ (sub_wire1[31] & 1'b1);
q[31] = (sub_wire1[30] & 1'b1) ^ (sub_wire1[31] & 1'b1) ^ (sub_wire1[0] & 1'b1);
    end
	 
end
	
	dcfifo_mixed_widths	dcfifo_mixed_widths_component (
				.rdclk (rdclk),
				.wrclk (wrclk),
				.wrreq (wrreq),
				.aclr (aclr),
				.data (data),
				.rdreq (rdreq),
				.wrfull (sub_wire0),
				.q (sub_wire1),
				.rdempty (sub_wire2),
				.wrusedw (sub_wire3),
				.rdusedw (sub_wire4),
				.rdfull (),
				.wrempty ());
	defparam
		dcfifo_mixed_widths_component.intended_device_family = "Cyclone IV E",
		dcfifo_mixed_widths_component.lpm_numwords = 4096,
		dcfifo_mixed_widths_component.lpm_showahead = "OFF",
		dcfifo_mixed_widths_component.lpm_type = "dcfifo_mixed_widths",
		dcfifo_mixed_widths_component.lpm_width = 8,
		dcfifo_mixed_widths_component.lpm_widthu = 12,
		dcfifo_mixed_widths_component.lpm_widthu_r = 10,
		dcfifo_mixed_widths_component.lpm_width_r = 32,
		dcfifo_mixed_widths_component.overflow_checking = "ON",
		dcfifo_mixed_widths_component.rdsync_delaypipe = 4,
		dcfifo_mixed_widths_component.read_aclr_synch = "OFF",
		dcfifo_mixed_widths_component.underflow_checking = "ON",
		dcfifo_mixed_widths_component.use_eab = "ON",
		dcfifo_mixed_widths_component.write_aclr_synch = "OFF",
		dcfifo_mixed_widths_component.wrsync_delaypipe = 4;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: AlmostEmpty NUMERIC "0"
// Retrieval info: PRIVATE: AlmostEmptyThr NUMERIC "-1"
// Retrieval info: PRIVATE: AlmostFull NUMERIC "0"
// Retrieval info: PRIVATE: AlmostFullThr NUMERIC "-1"
// Retrieval info: PRIVATE: CLOCKS_ARE_SYNCHRONIZED NUMERIC "0"
// Retrieval info: PRIVATE: Clock NUMERIC "4"
// Retrieval info: PRIVATE: Depth NUMERIC "4096"
// Retrieval info: PRIVATE: Empty NUMERIC "1"
// Retrieval info: PRIVATE: Full NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: LE_BasedFIFO NUMERIC "0"
// Retrieval info: PRIVATE: LegacyRREQ NUMERIC "1"
// Retrieval info: PRIVATE: MAX_DEPTH_BY_9 NUMERIC "0"
// Retrieval info: PRIVATE: OVERFLOW_CHECKING NUMERIC "0"
// Retrieval info: PRIVATE: Optimize NUMERIC "0"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: UNDERFLOW_CHECKING NUMERIC "0"
// Retrieval info: PRIVATE: UsedW NUMERIC "1"
// Retrieval info: PRIVATE: Width NUMERIC "8"
// Retrieval info: PRIVATE: dc_aclr NUMERIC "1"
// Retrieval info: PRIVATE: diff_widths NUMERIC "1"
// Retrieval info: PRIVATE: msb_usedw NUMERIC "0"
// Retrieval info: PRIVATE: output_width NUMERIC "32"
// Retrieval info: PRIVATE: rsEmpty NUMERIC "1"
// Retrieval info: PRIVATE: rsFull NUMERIC "0"
// Retrieval info: PRIVATE: rsUsedW NUMERIC "1"
// Retrieval info: PRIVATE: sc_aclr NUMERIC "0"
// Retrieval info: PRIVATE: sc_sclr NUMERIC "0"
// Retrieval info: PRIVATE: wsEmpty NUMERIC "0"
// Retrieval info: PRIVATE: wsFull NUMERIC "1"
// Retrieval info: PRIVATE: wsUsedW NUMERIC "1"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: CONSTANT: LPM_NUMWORDS NUMERIC "4096"
// Retrieval info: CONSTANT: LPM_SHOWAHEAD STRING "OFF"
// Retrieval info: CONSTANT: LPM_TYPE STRING "dcfifo_mixed_widths"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "8"
// Retrieval info: CONSTANT: LPM_WIDTHU NUMERIC "12"
// Retrieval info: CONSTANT: LPM_WIDTHU_R NUMERIC "10"
// Retrieval info: CONSTANT: LPM_WIDTH_R NUMERIC "32"
// Retrieval info: CONSTANT: OVERFLOW_CHECKING STRING "ON"
// Retrieval info: CONSTANT: RDSYNC_DELAYPIPE NUMERIC "4"
// Retrieval info: CONSTANT: READ_ACLR_SYNCH STRING "OFF"
// Retrieval info: CONSTANT: UNDERFLOW_CHECKING STRING "ON"
// Retrieval info: CONSTANT: USE_EAB STRING "ON"
// Retrieval info: CONSTANT: WRITE_ACLR_SYNCH STRING "OFF"
// Retrieval info: CONSTANT: WRSYNC_DELAYPIPE NUMERIC "4"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT GND "aclr"
// Retrieval info: USED_PORT: data 0 0 8 0 INPUT NODEFVAL "data[7..0]"
// Retrieval info: USED_PORT: q 0 0 32 0 OUTPUT NODEFVAL "q[31..0]"
// Retrieval info: USED_PORT: rdclk 0 0 0 0 INPUT NODEFVAL "rdclk"
// Retrieval info: USED_PORT: rdempty 0 0 0 0 OUTPUT NODEFVAL "rdempty"
// Retrieval info: USED_PORT: rdreq 0 0 0 0 INPUT NODEFVAL "rdreq"
// Retrieval info: USED_PORT: rdusedw 0 0 10 0 OUTPUT NODEFVAL "rdusedw[9..0]"
// Retrieval info: USED_PORT: wrclk 0 0 0 0 INPUT NODEFVAL "wrclk"
// Retrieval info: USED_PORT: wrfull 0 0 0 0 OUTPUT NODEFVAL "wrfull"
// Retrieval info: USED_PORT: wrreq 0 0 0 0 INPUT NODEFVAL "wrreq"
// Retrieval info: USED_PORT: wrusedw 0 0 12 0 OUTPUT NODEFVAL "wrusedw[11..0]"
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 8 0 data 0 0 8 0
// Retrieval info: CONNECT: @rdclk 0 0 0 0 rdclk 0 0 0 0
// Retrieval info: CONNECT: @rdreq 0 0 0 0 rdreq 0 0 0 0
// Retrieval info: CONNECT: @wrclk 0 0 0 0 wrclk 0 0 0 0
// Retrieval info: CONNECT: @wrreq 0 0 0 0 wrreq 0 0 0 0
// Retrieval info: CONNECT: q 0 0 32 0 @q 0 0 32 0
// Retrieval info: CONNECT: rdempty 0 0 0 0 @rdempty 0 0 0 0
// Retrieval info: CONNECT: rdusedw 0 0 10 0 @rdusedw 0 0 10 0
// Retrieval info: CONNECT: wrfull 0 0 0 0 @wrfull 0 0 0 0
// Retrieval info: CONNECT: wrusedw 0 0 12 0 @wrusedw 0 0 12 0
// Retrieval info: GEN_FILE: TYPE_NORMAL cmos1_fifo.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL cmos1_fifo.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL cmos1_fifo.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL cmos1_fifo.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL cmos1_fifo_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL cmos1_fifo_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
