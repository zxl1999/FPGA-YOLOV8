`timescale 1 ps/ 1 ps

module top_fpga(
	clk,
	rst_n,
	cam_scl,
	cam_sda,
	cam_data,
	cam_vsync,
	cam_hsync,
	cam_pclk,
	cam_xclk,
	cam_pdown,
	cam_reset,
	e_txen,
	e_tx,
	e_rxer,
	e_rxdv,
	e_rxclk,
	e_rx,
	led);
input	clk;
input	rst_n;
output	cam_scl;
inout	cam_sda;
input	[7:0] cam_data;
input	cam_vsync;
input	cam_hsync;
input	cam_pclk;
output	cam_xclk;
output	cam_pdown;
output	cam_reset;
output	e_txen;
output	[1:0] e_tx;
input	e_rxer;
input	e_rxdv;
input	e_rxclk;
input	[1:0] e_rx;
output	led;

//wire	gnd;
//wire	vcc;
wire	\Add0~0_combout ;
wire	\Add0~1 ;
wire	\Add0~2_combout ;
wire	\Add0~3 ;
wire	\Add0~4_combout ;
wire	\Add0~5 ;
wire	\Add0~6_combout ;
wire	\Add0~7 ;
wire	\Add0~8_combout ;
wire	AsyncReset_X11_Y15_GND;
wire	AsyncReset_X12_Y12_GND;
wire	AsyncReset_X12_Y14_GND;
wire	AsyncReset_X12_Y15_GND;
wire	AsyncReset_X1_Y17_GND;
wire	AsyncReset_X1_Y7_GND;
wire	AsyncReset_X24_Y15_GND;
wire	AsyncReset_X28_Y14_GND;
wire	AsyncReset_X28_Y15_GND;
wire	AsyncReset_X28_Y18_GND;
wire	AsyncReset_X2_Y7_GND;
wire	AsyncReset_X4_Y7_GND;
wire	\Equal0~0_combout ;
wire	\Equal0~1_combout ;
wire	\Equal0~2_combout ;
wire	\Equal0~3_combout ;
wire	\Equal0~4_combout ;
wire	\Equal0~5_combout ;
wire	\Equal0~6_combout ;
wire	\Equal0~7_combout ;
wire	\LessThan0~0_combout ;
wire	SyncLoad_X12_Y13_VCC;
wire	SyncLoad_X12_Y14_GND;
wire	SyncLoad_X12_Y15_GND;
wire	SyncLoad_X13_Y12_VCC;
wire	SyncLoad_X14_Y12_VCC;
wire	SyncLoad_X14_Y13_VCC;
wire	SyncLoad_X14_Y17_GND;
wire	SyncLoad_X16_Y11_VCC;
wire	SyncLoad_X16_Y12_VCC;
wire	SyncLoad_X16_Y13_VCC;
wire	SyncLoad_X17_Y13_VCC;
wire	SyncLoad_X1_Y17_GND;
wire	SyncLoad_X1_Y7_VCC;
wire	SyncLoad_X22_Y16_GND;
wire	SyncLoad_X22_Y19_VCC;
wire	SyncLoad_X22_Y8_VCC;
wire	SyncLoad_X23_Y15_GND;
wire	SyncLoad_X23_Y16_VCC;
wire	SyncLoad_X23_Y18_VCC;
wire	SyncLoad_X23_Y19_VCC;
wire	SyncLoad_X23_Y8_GND;
wire	SyncLoad_X24_Y16_GND;
wire	SyncLoad_X2_Y7_GND;
wire	SyncLoad_X4_Y7_VCC;
wire	SyncReset_X12_Y13_GND;
wire	SyncReset_X13_Y12_GND;
wire	SyncReset_X14_Y12_GND;
wire	SyncReset_X14_Y13_GND;
wire	SyncReset_X16_Y11_GND;
wire	SyncReset_X16_Y12_GND;
wire	SyncReset_X16_Y13_GND;
wire	SyncReset_X17_Y13_GND;
wire	SyncReset_X1_Y7_GND;
wire	SyncReset_X22_Y19_GND;
wire	SyncReset_X22_Y8_GND;
wire	SyncReset_X23_Y16_GND;
wire	SyncReset_X23_Y18_GND;
wire	SyncReset_X23_Y19_GND;
wire	SyncReset_X28_Y14_GND;
wire	SyncReset_X28_Y15_GND;
wire	SyncReset_X4_Y7_GND;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X14_Y17_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y16_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y17_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y18_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y17_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y17_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X19_Y12_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y19_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y16_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y8_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y18_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y19_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y16_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y14_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y15_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y15_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~combout ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ;
wire	[4:0] \alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus ;
//wire	\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [0];
//wire	\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [1];
//wire	\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [2];
//wire	\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [3];
//wire	\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [4];
wire	\alt_pll_inst|altpll_component|auto_generated|pll_lock_sync~feeder_combout ;
wire	\alt_pll_inst|altpll_component|auto_generated|pll_lock_sync~q ;
wire	[4:0] \alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk ;
//wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk [0];
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X17_Y17_SIG_VCC ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X22_Y8_SIG_VCC ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X18_Y17_SIG_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y16_SIG_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y17_SIG_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y18_SIG_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y17_SIG_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y17_SIG_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X14_Y17_SIG_SIG ;
//wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk [1];
//wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk [2];
//wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk [3];
//wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk [4];
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_fbout ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked_X17_Y1_SIG_VCC ;
wire	\cam_data[0]~input_o ;
wire	\cam_data[1]~input_o ;
wire	\cam_data[2]~input_o ;
wire	\cam_data[3]~input_o ;
wire	\cam_data[4]~input_o ;
wire	\cam_data[5]~input_o ;
wire	\cam_data[6]~input_o ;
wire	\cam_data[7]~input_o ;
wire	\cam_hsync~input_o ;
wire	\cam_pclk~input_o ;
wire	\cam_pclk~input_o_X12_Y13_SIG_VCC ;
wire	\cam_pclk~input_o_X13_Y12_SIG_VCC ;
wire	\cam_pclk~input_o_X13_Y13_SIG_VCC ;
wire	\cam_pclk~input_o_X14_Y13_SIG_VCC ;
wire	\cam_pclk~input_o_X16_Y13_SIG_VCC ;
wire	\cam_pclk~input_o_X17_Y13_SIG_VCC ;
wire	\cam_pclk~input_o_X1_Y7_SIG_VCC ;
wire	\cam_pclk~input_o_X2_Y7_SIG_VCC ;
wire	\cam_pclk~input_o_X3_Y7_SIG_VCC ;
wire	\cam_pclk~input_o_X4_Y7_SIG_VCC ;
wire	\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ;
wire	\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X13_Y13_SIG_SIG ;
wire	\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y13_SIG_SIG ;
wire	\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y13_SIG_SIG ;
wire	\cam_sda~input_o ;
wire	\cam_vsync~input_o ;
wire	\camera_if_inst|Equal0~0_combout ;
wire	\camera_if_inst|Equal0~1_combout ;
wire	\camera_if_inst|Equal0~2_combout ;
wire	\camera_if_inst|Equal0~3_combout ;
wire	\camera_if_inst|Equal0~4_combout ;
wire	\camera_if_inst|Equal1~0_combout ;
wire	\camera_if_inst|Equal1~1_combout ;
wire	\camera_if_inst|Equal2~0_combout ;
wire	\camera_if_inst|Equal3~0_combout ;
wire	\camera_if_inst|Equal3~1_combout ;
wire	\camera_if_inst|Equal3~2_combout ;
wire	\camera_if_inst|Equal3~3_combout ;
wire	\camera_if_inst|Equal3~4_combout ;
wire	\camera_if_inst|Equal4~0_combout ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y13_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y12_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y12_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y14_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X3_Y7_SIG ;
wire	[7:0] \camera_if_inst|cam_data_r0 ;
//wire	\camera_if_inst|cam_data_r0 [0];
wire	\camera_if_inst|cam_data_r0[0]~feeder_combout ;
//wire	\camera_if_inst|cam_data_r0 [1];
//wire	\camera_if_inst|cam_data_r0 [2];
//wire	\camera_if_inst|cam_data_r0 [3];
//wire	\camera_if_inst|cam_data_r0 [4];
//wire	\camera_if_inst|cam_data_r0 [5];
wire	\camera_if_inst|cam_data_r0[5]~feeder_combout ;
//wire	\camera_if_inst|cam_data_r0 [6];
//wire	\camera_if_inst|cam_data_r0 [7];
wire	[7:0] \camera_if_inst|cam_data_r1 ;
//wire	\camera_if_inst|cam_data_r1 [0];
//wire	\camera_if_inst|cam_data_r1 [1];
//wire	\camera_if_inst|cam_data_r1 [2];
//wire	\camera_if_inst|cam_data_r1 [3];
//wire	\camera_if_inst|cam_data_r1 [4];
//wire	\camera_if_inst|cam_data_r1 [5];
//wire	\camera_if_inst|cam_data_r1 [6];
//wire	\camera_if_inst|cam_data_r1 [7];
wire	\camera_if_inst|cam_data_r1~0_combout ;
wire	\camera_if_inst|cam_data_r1~1_combout ;
wire	\camera_if_inst|cam_data_r1~2_combout ;
wire	\camera_if_inst|cam_data_r1~3_combout ;
wire	\camera_if_inst|cam_data_r1~4_combout ;
wire	\camera_if_inst|cam_data_r1~5_combout ;
wire	\camera_if_inst|cam_data_r1~6_combout ;
wire	\camera_if_inst|cam_data_r1~7_combout ;
wire	[4:0] \camera_if_inst|cam_hsync_r ;
//wire	\camera_if_inst|cam_hsync_r [0];
wire	\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ;
//wire	\camera_if_inst|cam_hsync_r [1];
//wire	\camera_if_inst|cam_hsync_r [2];
//wire	\camera_if_inst|cam_hsync_r [3];
//wire	\camera_if_inst|cam_hsync_r [4];
wire	\camera_if_inst|cam_hsync_r~0_combout ;
wire	\camera_if_inst|cam_hsync_r~1_combout ;
wire	[4:0] \camera_if_inst|cam_vsync_r ;
//wire	\camera_if_inst|cam_vsync_r [0];
wire	\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ;
//wire	\camera_if_inst|cam_vsync_r [1];
//wire	\camera_if_inst|cam_vsync_r [2];
//wire	\camera_if_inst|cam_vsync_r [3];
//wire	\camera_if_inst|cam_vsync_r [4];
wire	[3:0] \camera_if_inst|f_cnt ;
//wire	\camera_if_inst|f_cnt [0];
wire	\camera_if_inst|f_cnt[0]~5_combout ;
//wire	\camera_if_inst|f_cnt [1];
wire	\camera_if_inst|f_cnt[1]~4_combout ;
//wire	\camera_if_inst|f_cnt [2];
wire	\camera_if_inst|f_cnt[2]~3_combout ;
//wire	\camera_if_inst|f_cnt [3];
wire	\camera_if_inst|f_cnt[3]~2_combout ;
wire	\camera_if_inst|f_cnt[3]~6_combout ;
wire	[15:0] \camera_if_inst|h_cnt ;
//wire	\camera_if_inst|h_cnt [0];
wire	\camera_if_inst|h_cnt[0]~16_combout ;
wire	\camera_if_inst|h_cnt[0]~17 ;
//wire	\camera_if_inst|h_cnt [10];
wire	\camera_if_inst|h_cnt[10]~36_combout ;
wire	\camera_if_inst|h_cnt[10]~37 ;
//wire	\camera_if_inst|h_cnt [11];
wire	\camera_if_inst|h_cnt[11]~38_combout ;
wire	\camera_if_inst|h_cnt[11]~39 ;
//wire	\camera_if_inst|h_cnt [12];
wire	\camera_if_inst|h_cnt[12]~40_combout ;
wire	\camera_if_inst|h_cnt[12]~41 ;
//wire	\camera_if_inst|h_cnt [13];
wire	\camera_if_inst|h_cnt[13]~42_combout ;
wire	\camera_if_inst|h_cnt[13]~43 ;
//wire	\camera_if_inst|h_cnt [14];
wire	\camera_if_inst|h_cnt[14]~44_combout ;
wire	\camera_if_inst|h_cnt[14]~45 ;
//wire	\camera_if_inst|h_cnt [15];
wire	\camera_if_inst|h_cnt[15]~46_combout ;
//wire	\camera_if_inst|h_cnt [1];
wire	\camera_if_inst|h_cnt[1]~18_combout ;
wire	\camera_if_inst|h_cnt[1]~19 ;
//wire	\camera_if_inst|h_cnt [2];
wire	\camera_if_inst|h_cnt[2]~20_combout ;
wire	\camera_if_inst|h_cnt[2]~21 ;
//wire	\camera_if_inst|h_cnt [3];
wire	\camera_if_inst|h_cnt[3]~22_combout ;
wire	\camera_if_inst|h_cnt[3]~23 ;
//wire	\camera_if_inst|h_cnt [4];
wire	\camera_if_inst|h_cnt[4]~24_combout ;
wire	\camera_if_inst|h_cnt[4]~25 ;
//wire	\camera_if_inst|h_cnt [5];
wire	\camera_if_inst|h_cnt[5]~26_combout ;
wire	\camera_if_inst|h_cnt[5]~27 ;
//wire	\camera_if_inst|h_cnt [6];
wire	\camera_if_inst|h_cnt[6]~28_combout ;
wire	\camera_if_inst|h_cnt[6]~29 ;
//wire	\camera_if_inst|h_cnt [7];
wire	\camera_if_inst|h_cnt[7]~30_combout ;
wire	\camera_if_inst|h_cnt[7]~31 ;
//wire	\camera_if_inst|h_cnt [8];
wire	\camera_if_inst|h_cnt[8]~32_combout ;
wire	\camera_if_inst|h_cnt[8]~33 ;
//wire	\camera_if_inst|h_cnt [9];
wire	\camera_if_inst|h_cnt[9]~34_combout ;
wire	\camera_if_inst|h_cnt[9]~35 ;
wire	[7:0] \camera_if_inst|u_I2C_AV_Config|LUT_INDEX ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0]~22_combout ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1]~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1]~8 ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2]~10 ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2]~9_combout ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3]~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3]~12 ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4]~14_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4]~15 ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5]~16_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5]~17 ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6]~18_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6]~19 ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~20_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan0~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan0~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan0~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan0~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan1~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|Selector3~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|Selector3~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|Selector3~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~feeder_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~q ;
wire	\camera_if_inst|u_I2C_AV_Config|i2c_en_r1~q ;
wire	\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ;
wire	[15:0] \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [0];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0]~16_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0]~17 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [10];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10]~36_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10]~37 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [11];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11]~38_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11]~39 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [12];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12]~40_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12]~41 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [13];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13]~42_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13]~43 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [14];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14]~44_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14]~45 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [15];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15]~46_combout ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [1];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1]~18_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1]~19 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [2];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2]~20_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2]~21 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [3];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3]~22_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3]~23 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [4];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4]~24_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4]~25 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [5];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5]~26_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5]~27 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [6];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6]~28_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6]~29 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [7];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7]~30_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7]~31 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [8];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8]~32_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8]~33 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [9];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9]~34_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9]~35 ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~q ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X14_Y17_INV ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_GO~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_WR~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST.00~q ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST.10~q ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST~12_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST~13_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACK~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACK~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACK~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Equal0~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Equal0~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Equal3~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Equal3~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Equal5~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~12_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~13_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~14_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~15_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~16_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~17_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~18_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~19_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~20_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~21_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~22_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~23_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~24_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~25_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~26_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~27_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~28_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~29_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~30_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~31_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SDO~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SDO~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SDO~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SDO~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SDO~4_combout ;
wire	[5:0] \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER ;
//wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0];
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0]~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0]~7 ;
//wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1];
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1]~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1]~9 ;
//wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2];
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2]~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2]~11 ;
//wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3];
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3]~13_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3]~14 ;
//wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4];
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4]~15_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4]~16 ;
//wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5];
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~17_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector2~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector8~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector9~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector9~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|comb~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|comb~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9_combout ;
wire	[15:0] \camera_if_inst|v_cnt ;
//wire	\camera_if_inst|v_cnt [0];
wire	\camera_if_inst|v_cnt[0]~16_combout ;
wire	\camera_if_inst|v_cnt[0]~17 ;
//wire	\camera_if_inst|v_cnt [10];
wire	\camera_if_inst|v_cnt[10]~37_combout ;
wire	\camera_if_inst|v_cnt[10]~38 ;
//wire	\camera_if_inst|v_cnt [11];
wire	\camera_if_inst|v_cnt[11]~39_combout ;
wire	\camera_if_inst|v_cnt[11]~40 ;
//wire	\camera_if_inst|v_cnt [12];
wire	\camera_if_inst|v_cnt[12]~41_combout ;
wire	\camera_if_inst|v_cnt[12]~42 ;
//wire	\camera_if_inst|v_cnt [13];
wire	\camera_if_inst|v_cnt[13]~43_combout ;
wire	\camera_if_inst|v_cnt[13]~44 ;
//wire	\camera_if_inst|v_cnt [14];
wire	\camera_if_inst|v_cnt[14]~45_combout ;
wire	\camera_if_inst|v_cnt[14]~46 ;
//wire	\camera_if_inst|v_cnt [15];
wire	\camera_if_inst|v_cnt[15]~47_combout ;
//wire	\camera_if_inst|v_cnt [1];
wire	\camera_if_inst|v_cnt[1]~19_combout ;
wire	\camera_if_inst|v_cnt[1]~20 ;
//wire	\camera_if_inst|v_cnt [2];
wire	\camera_if_inst|v_cnt[2]~21_combout ;
wire	\camera_if_inst|v_cnt[2]~22 ;
//wire	\camera_if_inst|v_cnt [3];
wire	\camera_if_inst|v_cnt[3]~23_combout ;
wire	\camera_if_inst|v_cnt[3]~24 ;
//wire	\camera_if_inst|v_cnt [4];
wire	\camera_if_inst|v_cnt[4]~25_combout ;
wire	\camera_if_inst|v_cnt[4]~26 ;
//wire	\camera_if_inst|v_cnt [5];
wire	\camera_if_inst|v_cnt[5]~27_combout ;
wire	\camera_if_inst|v_cnt[5]~28 ;
//wire	\camera_if_inst|v_cnt [6];
wire	\camera_if_inst|v_cnt[6]~29_combout ;
wire	\camera_if_inst|v_cnt[6]~30 ;
//wire	\camera_if_inst|v_cnt [7];
wire	\camera_if_inst|v_cnt[7]~31_combout ;
wire	\camera_if_inst|v_cnt[7]~32 ;
//wire	\camera_if_inst|v_cnt [8];
wire	\camera_if_inst|v_cnt[8]~18_combout ;
wire	\camera_if_inst|v_cnt[8]~33_combout ;
wire	\camera_if_inst|v_cnt[8]~34 ;
//wire	\camera_if_inst|v_cnt [9];
wire	\camera_if_inst|v_cnt[9]~35_combout ;
wire	\camera_if_inst|v_cnt[9]~36 ;
wire	\clk_25m~0_combout ;
wire	\clk_25m~clkctrl_outclk ;
wire	\clk_25m~clkctrl_outclk_X12_Y13_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X13_Y12_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X14_Y12_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X16_Y11_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X17_Y12_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X17_Y13_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X17_Y14_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X22_Y19_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X23_Y16_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X23_Y18_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X24_Y15_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X25_Y16_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X3_Y7_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y12_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y11_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y12_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y19_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X22_Y19_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y14_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y15_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[3]~13_combout_X24_Y16_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X22_Y16_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout_X19_Y12_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y14_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y15_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y18_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y16_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y18_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X24_Y15_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X25_Y16_SIG_SIG ;
wire	\clk_25m~q ;
wire	\clk~input_o ;
wire	\clk~inputclkctrl_outclk ;
wire	\clk~inputclkctrl_outclk_X11_Y15_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X12_Y12_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ;
wire	\clk~inputclkctrl_outclk__reset_init[5]_X12_Y12_SIG_INV ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita0~COUT ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita0~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~COUT ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~combout ;
wire	[1:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [1];
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [0];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [10];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [2];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [3];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [4];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [5];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [6];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9]~feeder_combout ;
wire	[31:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [18];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [19];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [20];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [21];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [22];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [23];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [24];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [25];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [26];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [27];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [28];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [29];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [30];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [31];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [9];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [9];
wire	[7:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [7];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [9];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [8];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [9];
wire	[7:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [7];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [9];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [8];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [9];
wire	[7:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [7];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [9];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [8];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [9];
wire	[7:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3_PORTBDATAOUT_bus ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3_PORTBDATAOUT_bus [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3_PORTBDATAOUT_bus [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3_PORTBDATAOUT_bus [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3_PORTBDATAOUT_bus [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3_PORTBDATAOUT_bus [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3_PORTBDATAOUT_bus [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3_PORTBDATAOUT_bus [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3_PORTBDATAOUT_bus [7];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [9];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [8];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11_cout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~13 ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~15 ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~17 ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1_cout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3_cout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5_cout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7_cout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9_cout ;
wire	[11:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~1_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~2_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~3_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~5_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|data_wire[2]~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~10_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~1_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~7_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~8_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~9_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ;
wire	[2:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [2];
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [0];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0]~0_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [1];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [7];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor0~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor1~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor2~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor3~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor4~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor5~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor6~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor7~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor8~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor9~combout ;
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [9];
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor0~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor1~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor2~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor3~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor4~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor5~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor6~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor7~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor8~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor9~combout ;
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [0];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [10];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [1];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [2];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [3];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [4];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [5];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [6];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [7];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [8];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9]~feeder_combout ;
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [7];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9]~feeder_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~1_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~2_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~3_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~5_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|data_wire[2]~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~10_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~6_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~7_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~8_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~9_combout ;
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [10];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10]~0_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1]~8_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2]~7_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3]~9_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4]~5_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5]~6_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6]~3_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7]~4_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8]~1_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9]~2_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2~q ;
wire	[12:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0]~0_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [12];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9];
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [0];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [10];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [3];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [6];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9]~feeder_combout ;
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [10];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [3];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [5];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [7];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9]~feeder_combout ;
tri1	devclrn;
tri1	devoe;
tri1	devpor;
wire	\e_rx[0]~input_o ;
wire	\e_rx[1]~input_o ;
wire	\e_rxclk~input_o ;
wire	\e_rxclk~input_o_X23_Y19_INV_VCC ;
wire	\e_rxclk~input_o_X33_Y15_INV_VCC ;
wire	\e_rxclk~input_o__mii_to_rmii_inst|tx_dv_reg~q_X23_Y19_SIG_SIG ;
wire	\e_rxdv~input_o ;
wire	\e_rxer~input_o ;
wire	[31:0] \eth_udp_inst|crc32_inst|crc_data ;
//wire	\eth_udp_inst|crc32_inst|crc_data [0];
//wire	\eth_udp_inst|crc32_inst|crc_data [10];
//wire	\eth_udp_inst|crc32_inst|crc_data [11];
//wire	\eth_udp_inst|crc32_inst|crc_data [12];
//wire	\eth_udp_inst|crc32_inst|crc_data [13];
//wire	\eth_udp_inst|crc32_inst|crc_data [14];
//wire	\eth_udp_inst|crc32_inst|crc_data [15];
//wire	\eth_udp_inst|crc32_inst|crc_data [16];
//wire	\eth_udp_inst|crc32_inst|crc_data [17];
//wire	\eth_udp_inst|crc32_inst|crc_data [18];
//wire	\eth_udp_inst|crc32_inst|crc_data [19];
//wire	\eth_udp_inst|crc32_inst|crc_data [1];
//wire	\eth_udp_inst|crc32_inst|crc_data [20];
//wire	\eth_udp_inst|crc32_inst|crc_data [21];
//wire	\eth_udp_inst|crc32_inst|crc_data [22];
//wire	\eth_udp_inst|crc32_inst|crc_data [23];
//wire	\eth_udp_inst|crc32_inst|crc_data [24];
//wire	\eth_udp_inst|crc32_inst|crc_data [25];
//wire	\eth_udp_inst|crc32_inst|crc_data [26];
//wire	\eth_udp_inst|crc32_inst|crc_data [27];
//wire	\eth_udp_inst|crc32_inst|crc_data [28];
wire	\eth_udp_inst|crc32_inst|crc_data[28]~9_combout ;
//wire	\eth_udp_inst|crc32_inst|crc_data [29];
//wire	\eth_udp_inst|crc32_inst|crc_data [2];
//wire	\eth_udp_inst|crc32_inst|crc_data [30];
//wire	\eth_udp_inst|crc32_inst|crc_data [31];
//wire	\eth_udp_inst|crc32_inst|crc_data [3];
//wire	\eth_udp_inst|crc32_inst|crc_data [4];
//wire	\eth_udp_inst|crc32_inst|crc_data [5];
//wire	\eth_udp_inst|crc32_inst|crc_data [6];
//wire	\eth_udp_inst|crc32_inst|crc_data [7];
//wire	\eth_udp_inst|crc32_inst|crc_data [8];
//wire	\eth_udp_inst|crc32_inst|crc_data [9];
wire	\eth_udp_inst|crc32_inst|crc_data~10_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~11_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~12_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~13_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~14_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~15_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~16_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~17_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~18_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~19_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~20_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~21_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~22_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~23_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~24_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~25_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~26_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~27_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~28_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~29_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~30_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~31_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~32_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~33_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~34_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~35_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~36_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~37_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~38_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~39_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~40_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~8_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next[28]~1_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next[29]~0_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next~2_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next~3_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next~4_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next~5_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next~6_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next~7_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~1 ;
wire	\eth_udp_inst|ip_send_inst|Add13~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~11 ;
wire	\eth_udp_inst|ip_send_inst|Add13~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~13 ;
wire	\eth_udp_inst|ip_send_inst|Add13~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~15 ;
wire	\eth_udp_inst|ip_send_inst|Add13~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~17 ;
wire	\eth_udp_inst|ip_send_inst|Add13~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~19 ;
wire	\eth_udp_inst|ip_send_inst|Add13~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~21 ;
wire	\eth_udp_inst|ip_send_inst|Add13~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~23 ;
wire	\eth_udp_inst|ip_send_inst|Add13~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~25 ;
wire	\eth_udp_inst|ip_send_inst|Add13~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~27 ;
wire	\eth_udp_inst|ip_send_inst|Add13~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~29 ;
wire	\eth_udp_inst|ip_send_inst|Add13~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~3 ;
wire	\eth_udp_inst|ip_send_inst|Add13~30_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~5 ;
wire	\eth_udp_inst|ip_send_inst|Add13~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~7 ;
wire	\eth_udp_inst|ip_send_inst|Add13~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~9 ;
wire	\eth_udp_inst|ip_send_inst|Add2~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~1 ;
wire	\eth_udp_inst|ip_send_inst|Add2~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~11 ;
wire	\eth_udp_inst|ip_send_inst|Add2~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~13 ;
wire	\eth_udp_inst|ip_send_inst|Add2~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~15 ;
wire	\eth_udp_inst|ip_send_inst|Add2~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~17 ;
wire	\eth_udp_inst|ip_send_inst|Add2~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~19 ;
wire	\eth_udp_inst|ip_send_inst|Add2~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~21 ;
wire	\eth_udp_inst|ip_send_inst|Add2~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~23 ;
wire	\eth_udp_inst|ip_send_inst|Add2~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~25 ;
wire	\eth_udp_inst|ip_send_inst|Add2~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~27 ;
wire	\eth_udp_inst|ip_send_inst|Add2~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~3 ;
wire	\eth_udp_inst|ip_send_inst|Add2~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~5 ;
wire	\eth_udp_inst|ip_send_inst|Add2~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~7 ;
wire	\eth_udp_inst|ip_send_inst|Add2~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~9 ;
wire	\eth_udp_inst|ip_send_inst|Add3~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add3~1 ;
wire	\eth_udp_inst|ip_send_inst|Add3~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add3~3 ;
wire	\eth_udp_inst|ip_send_inst|Add3~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~1 ;
wire	\eth_udp_inst|ip_send_inst|Add4~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~11 ;
wire	\eth_udp_inst|ip_send_inst|Add4~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~13 ;
wire	\eth_udp_inst|ip_send_inst|Add4~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~15 ;
wire	\eth_udp_inst|ip_send_inst|Add4~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~17 ;
wire	\eth_udp_inst|ip_send_inst|Add4~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~19 ;
wire	\eth_udp_inst|ip_send_inst|Add4~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~21 ;
wire	\eth_udp_inst|ip_send_inst|Add4~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~23 ;
wire	\eth_udp_inst|ip_send_inst|Add4~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~25 ;
wire	\eth_udp_inst|ip_send_inst|Add4~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~27 ;
wire	\eth_udp_inst|ip_send_inst|Add4~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~29 ;
wire	\eth_udp_inst|ip_send_inst|Add4~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~3 ;
wire	\eth_udp_inst|ip_send_inst|Add4~30_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~31 ;
wire	\eth_udp_inst|ip_send_inst|Add4~32_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~33 ;
wire	\eth_udp_inst|ip_send_inst|Add4~34_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~5 ;
wire	\eth_udp_inst|ip_send_inst|Add4~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~7 ;
wire	\eth_udp_inst|ip_send_inst|Add4~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~9 ;
wire	\eth_udp_inst|ip_send_inst|Add5~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~1 ;
wire	\eth_udp_inst|ip_send_inst|Add5~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~11 ;
wire	\eth_udp_inst|ip_send_inst|Add5~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~13 ;
wire	\eth_udp_inst|ip_send_inst|Add5~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~15 ;
wire	\eth_udp_inst|ip_send_inst|Add5~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~17 ;
wire	\eth_udp_inst|ip_send_inst|Add5~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~19 ;
wire	\eth_udp_inst|ip_send_inst|Add5~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~21 ;
wire	\eth_udp_inst|ip_send_inst|Add5~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~23 ;
wire	\eth_udp_inst|ip_send_inst|Add5~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~25 ;
wire	\eth_udp_inst|ip_send_inst|Add5~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~27 ;
wire	\eth_udp_inst|ip_send_inst|Add5~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~29 ;
wire	\eth_udp_inst|ip_send_inst|Add5~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~3 ;
wire	\eth_udp_inst|ip_send_inst|Add5~30_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~31 ;
wire	\eth_udp_inst|ip_send_inst|Add5~32_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~33 ;
wire	\eth_udp_inst|ip_send_inst|Add5~34_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~5 ;
wire	\eth_udp_inst|ip_send_inst|Add5~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~7 ;
wire	\eth_udp_inst|ip_send_inst|Add5~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~9 ;
wire	\eth_udp_inst|ip_send_inst|Add6~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~1 ;
wire	\eth_udp_inst|ip_send_inst|Add6~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~11 ;
wire	\eth_udp_inst|ip_send_inst|Add6~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~13 ;
wire	\eth_udp_inst|ip_send_inst|Add6~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~15 ;
wire	\eth_udp_inst|ip_send_inst|Add6~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~17 ;
wire	\eth_udp_inst|ip_send_inst|Add6~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~19 ;
wire	\eth_udp_inst|ip_send_inst|Add6~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~21 ;
wire	\eth_udp_inst|ip_send_inst|Add6~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~23 ;
wire	\eth_udp_inst|ip_send_inst|Add6~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~25 ;
wire	\eth_udp_inst|ip_send_inst|Add6~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~27 ;
wire	\eth_udp_inst|ip_send_inst|Add6~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~3 ;
wire	\eth_udp_inst|ip_send_inst|Add6~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~5 ;
wire	\eth_udp_inst|ip_send_inst|Add6~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~7 ;
wire	\eth_udp_inst|ip_send_inst|Add6~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~9 ;
wire	\eth_udp_inst|ip_send_inst|Add7~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~1 ;
wire	\eth_udp_inst|ip_send_inst|Add7~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~11 ;
wire	\eth_udp_inst|ip_send_inst|Add7~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~13 ;
wire	\eth_udp_inst|ip_send_inst|Add7~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~15 ;
wire	\eth_udp_inst|ip_send_inst|Add7~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~17 ;
wire	\eth_udp_inst|ip_send_inst|Add7~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~19 ;
wire	\eth_udp_inst|ip_send_inst|Add7~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~21 ;
wire	\eth_udp_inst|ip_send_inst|Add7~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~23 ;
wire	\eth_udp_inst|ip_send_inst|Add7~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~25 ;
wire	\eth_udp_inst|ip_send_inst|Add7~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~27 ;
wire	\eth_udp_inst|ip_send_inst|Add7~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~29 ;
wire	\eth_udp_inst|ip_send_inst|Add7~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~3 ;
wire	\eth_udp_inst|ip_send_inst|Add7~30_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~31 ;
wire	\eth_udp_inst|ip_send_inst|Add7~32_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~5 ;
wire	\eth_udp_inst|ip_send_inst|Add7~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~7 ;
wire	\eth_udp_inst|ip_send_inst|Add7~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~9 ;
wire	\eth_udp_inst|ip_send_inst|Add8~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~1 ;
wire	\eth_udp_inst|ip_send_inst|Add8~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~11 ;
wire	\eth_udp_inst|ip_send_inst|Add8~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~13 ;
wire	\eth_udp_inst|ip_send_inst|Add8~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~15 ;
wire	\eth_udp_inst|ip_send_inst|Add8~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~17 ;
wire	\eth_udp_inst|ip_send_inst|Add8~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~19 ;
wire	\eth_udp_inst|ip_send_inst|Add8~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~21 ;
wire	\eth_udp_inst|ip_send_inst|Add8~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~23 ;
wire	\eth_udp_inst|ip_send_inst|Add8~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~25 ;
wire	\eth_udp_inst|ip_send_inst|Add8~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~27 ;
wire	\eth_udp_inst|ip_send_inst|Add8~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~29 ;
wire	\eth_udp_inst|ip_send_inst|Add8~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~3 ;
wire	\eth_udp_inst|ip_send_inst|Add8~30_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~5 ;
wire	\eth_udp_inst|ip_send_inst|Add8~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~7 ;
wire	\eth_udp_inst|ip_send_inst|Add8~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~9 ;
wire	\eth_udp_inst|ip_send_inst|Add9~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~1 ;
wire	\eth_udp_inst|ip_send_inst|Add9~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~11 ;
wire	\eth_udp_inst|ip_send_inst|Add9~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~13 ;
wire	\eth_udp_inst|ip_send_inst|Add9~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~15 ;
wire	\eth_udp_inst|ip_send_inst|Add9~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~17 ;
wire	\eth_udp_inst|ip_send_inst|Add9~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~19 ;
wire	\eth_udp_inst|ip_send_inst|Add9~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~21 ;
wire	\eth_udp_inst|ip_send_inst|Add9~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~23 ;
wire	\eth_udp_inst|ip_send_inst|Add9~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~25 ;
wire	\eth_udp_inst|ip_send_inst|Add9~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~27 ;
wire	\eth_udp_inst|ip_send_inst|Add9~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~29 ;
wire	\eth_udp_inst|ip_send_inst|Add9~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~3 ;
wire	\eth_udp_inst|ip_send_inst|Add9~30_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~31 ;
wire	\eth_udp_inst|ip_send_inst|Add9~32_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~33 ;
wire	\eth_udp_inst|ip_send_inst|Add9~34_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~35 ;
wire	\eth_udp_inst|ip_send_inst|Add9~36_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~5 ;
wire	\eth_udp_inst|ip_send_inst|Add9~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~7 ;
wire	\eth_udp_inst|ip_send_inst|Add9~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~9 ;
wire	\eth_udp_inst|ip_send_inst|Equal1~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal1~1_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y14_SIG ;
wire	\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y15_SIG ;
wire	\eth_udp_inst|ip_send_inst|Equal8~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal8~1_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal8~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal8~3_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal8~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal8~5_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal8~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal9~0_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~0_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~1_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~2_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~3_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~4_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~5_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~6_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~7_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan2~0_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan2~1_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan2~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux13~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux13~1_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux13~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux13~3_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux13~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux16~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux17~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux17~1_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux20~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux21~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux24~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux24~1_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux25~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux27~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux28~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux29~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux31~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux32~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux33~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux35~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux35~1_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux36~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux37~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux39~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux40~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux41~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux43~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux44~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux45~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux47~0_combout ;
wire	\eth_udp_inst|ip_send_inst|always10~0_combout ;
wire	\eth_udp_inst|ip_send_inst|always11~0_combout ;
wire	\eth_udp_inst|ip_send_inst|always13~0_combout ;
wire	\eth_udp_inst|ip_send_inst|always16~0_combout ;
wire	\eth_udp_inst|ip_send_inst|always3~2_combout ;
wire	\eth_udp_inst|ip_send_inst|always3~3_combout ;
wire	\eth_udp_inst|ip_send_inst|always3~4_combout ;
wire	\eth_udp_inst|ip_send_inst|always7~0_combout ;
wire	\eth_udp_inst|ip_send_inst|always7~1_combout ;
wire	[31:0] \eth_udp_inst|ip_send_inst|check_sum ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [0];
wire	\eth_udp_inst|ip_send_inst|check_sum[0]~17_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[0]~18 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [10];
wire	\eth_udp_inst|ip_send_inst|check_sum[10]~37_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[10]~38 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [11];
wire	\eth_udp_inst|ip_send_inst|check_sum[11]~39_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[11]~40 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [12];
wire	\eth_udp_inst|ip_send_inst|check_sum[12]~41_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[12]~42 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [13];
wire	\eth_udp_inst|ip_send_inst|check_sum[13]~43_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[13]~44 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [14];
wire	\eth_udp_inst|ip_send_inst|check_sum[14]~45_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[14]~46 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [15];
wire	\eth_udp_inst|ip_send_inst|check_sum[15]~48_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[15]~49 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [16];
wire	\eth_udp_inst|ip_send_inst|check_sum[16]~52_combout ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [17];
//wire	\eth_udp_inst|ip_send_inst|check_sum [18];
//wire	\eth_udp_inst|ip_send_inst|check_sum [19];
//wire	\eth_udp_inst|ip_send_inst|check_sum [1];
wire	\eth_udp_inst|ip_send_inst|check_sum[1]~19_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[1]~20 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [20];
//wire	\eth_udp_inst|ip_send_inst|check_sum [21];
//wire	\eth_udp_inst|ip_send_inst|check_sum [22];
//wire	\eth_udp_inst|ip_send_inst|check_sum [23];
//wire	\eth_udp_inst|ip_send_inst|check_sum [24];
//wire	\eth_udp_inst|ip_send_inst|check_sum [25];
//wire	\eth_udp_inst|ip_send_inst|check_sum [26];
//wire	\eth_udp_inst|ip_send_inst|check_sum [27];
//wire	\eth_udp_inst|ip_send_inst|check_sum [28];
//wire	\eth_udp_inst|ip_send_inst|check_sum [29];
//wire	\eth_udp_inst|ip_send_inst|check_sum [2];
wire	\eth_udp_inst|ip_send_inst|check_sum[2]~21_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[2]~22 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [30];
//wire	\eth_udp_inst|ip_send_inst|check_sum [31];
//wire	\eth_udp_inst|ip_send_inst|check_sum [3];
wire	\eth_udp_inst|ip_send_inst|check_sum[3]~23_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[3]~24 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [4];
wire	\eth_udp_inst|ip_send_inst|check_sum[4]~25_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[4]~26 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [5];
wire	\eth_udp_inst|ip_send_inst|check_sum[5]~27_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[5]~28 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [6];
wire	\eth_udp_inst|ip_send_inst|check_sum[6]~29_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[6]~30 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [7];
wire	\eth_udp_inst|ip_send_inst|check_sum[7]~31_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[7]~32 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [8];
wire	\eth_udp_inst|ip_send_inst|check_sum[8]~33_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[8]~34 ;
wire	\eth_udp_inst|ip_send_inst|check_sum[8]~47_combout ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [9];
wire	\eth_udp_inst|ip_send_inst|check_sum[9]~35_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[9]~36 ;
wire	\eth_udp_inst|ip_send_inst|check_sum~50_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum~51_combout ;
wire	[4:0] \eth_udp_inst|ip_send_inst|cnt ;
//wire	\eth_udp_inst|ip_send_inst|cnt [0];
wire	\eth_udp_inst|ip_send_inst|cnt[0]~5_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt[0]~6 ;
//wire	\eth_udp_inst|ip_send_inst|cnt [1];
wire	\eth_udp_inst|ip_send_inst|cnt[1]~7_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt[1]~8 ;
//wire	\eth_udp_inst|ip_send_inst|cnt [2];
wire	\eth_udp_inst|ip_send_inst|cnt[2]~10 ;
wire	\eth_udp_inst|ip_send_inst|cnt[2]~9_combout ;
//wire	\eth_udp_inst|ip_send_inst|cnt [3];
wire	\eth_udp_inst|ip_send_inst|cnt[3]~11_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt[3]~11_combout__SyncReset_X24_Y16_SIG ;
wire	\eth_udp_inst|ip_send_inst|cnt[3]~12_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt[3]~13_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt[3]~14_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt[3]~15 ;
//wire	\eth_udp_inst|ip_send_inst|cnt [4];
wire	\eth_udp_inst|ip_send_inst|cnt[4]~16_combout ;
wire	[4:0] \eth_udp_inst|ip_send_inst|cnt_add ;
//wire	\eth_udp_inst|ip_send_inst|cnt_add [0];
wire	\eth_udp_inst|ip_send_inst|cnt_add[0]~5_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_add[0]~6 ;
//wire	\eth_udp_inst|ip_send_inst|cnt_add [1];
wire	\eth_udp_inst|ip_send_inst|cnt_add[1]~7_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_add[1]~8 ;
//wire	\eth_udp_inst|ip_send_inst|cnt_add [2];
wire	\eth_udp_inst|ip_send_inst|cnt_add[2]~10 ;
wire	\eth_udp_inst|ip_send_inst|cnt_add[2]~9_combout ;
//wire	\eth_udp_inst|ip_send_inst|cnt_add [3];
wire	\eth_udp_inst|ip_send_inst|cnt_add[3]~11_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_add[3]~12 ;
//wire	\eth_udp_inst|ip_send_inst|cnt_add [4];
wire	\eth_udp_inst|ip_send_inst|cnt_add[4]~13_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_add[4]~15_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout ;
wire	[2:0] \eth_udp_inst|ip_send_inst|cnt_send_bit ;
//wire	\eth_udp_inst|ip_send_inst|cnt_send_bit [0];
//wire	\eth_udp_inst|ip_send_inst|cnt_send_bit [1];
//wire	\eth_udp_inst|ip_send_inst|cnt_send_bit [2];
wire	\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_send_bit~2_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_send_bit~4_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_send_bit~5_combout ;
wire	\eth_udp_inst|ip_send_inst|crc_clr~q ;
wire	\eth_udp_inst|ip_send_inst|crc_en~q ;
wire	[15:0] \eth_udp_inst|ip_send_inst|data_cnt ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [0];
wire	\eth_udp_inst|ip_send_inst|data_cnt[0]~16_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[0]~17 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [10];
wire	\eth_udp_inst|ip_send_inst|data_cnt[10]~36_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[10]~37 ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [11];
wire	\eth_udp_inst|ip_send_inst|data_cnt[11]~42_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[11]~43 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [12];
wire	\eth_udp_inst|ip_send_inst|data_cnt[12]~44_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[12]~45 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [13];
wire	\eth_udp_inst|ip_send_inst|data_cnt[13]~46_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[13]~47 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [14];
wire	\eth_udp_inst|ip_send_inst|data_cnt[14]~48_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[14]~49 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [15];
wire	\eth_udp_inst|ip_send_inst|data_cnt[15]~50_combout ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [1];
wire	\eth_udp_inst|ip_send_inst|data_cnt[1]~18_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[1]~19 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [2];
wire	\eth_udp_inst|ip_send_inst|data_cnt[2]~20_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[2]~21 ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[2]~38_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[2]~39_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[2]~40_combout ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [3];
wire	\eth_udp_inst|ip_send_inst|data_cnt[3]~22_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[3]~23 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [4];
wire	\eth_udp_inst|ip_send_inst|data_cnt[4]~24_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[4]~25 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [5];
wire	\eth_udp_inst|ip_send_inst|data_cnt[5]~26_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[5]~27 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [6];
wire	\eth_udp_inst|ip_send_inst|data_cnt[6]~28_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[6]~29 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [7];
wire	\eth_udp_inst|ip_send_inst|data_cnt[7]~30_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[7]~31 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [8];
wire	\eth_udp_inst|ip_send_inst|data_cnt[8]~32_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[8]~33 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [9];
wire	\eth_udp_inst|ip_send_inst|data_cnt[9]~34_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[9]~35 ;
wire	[15:0] \eth_udp_inst|ip_send_inst|data_len ;
//wire	\eth_udp_inst|ip_send_inst|data_len [0];
//wire	\eth_udp_inst|ip_send_inst|data_len [10];
wire	\eth_udp_inst|ip_send_inst|data_len[10]~0_combout ;
//wire	\eth_udp_inst|ip_send_inst|data_len [11];
//wire	\eth_udp_inst|ip_send_inst|data_len [12];
//wire	\eth_udp_inst|ip_send_inst|data_len [13];
//wire	\eth_udp_inst|ip_send_inst|data_len [14];
//wire	\eth_udp_inst|ip_send_inst|data_len [15];
//wire	\eth_udp_inst|ip_send_inst|data_len [1];
//wire	\eth_udp_inst|ip_send_inst|data_len [2];
//wire	\eth_udp_inst|ip_send_inst|data_len [3];
//wire	\eth_udp_inst|ip_send_inst|data_len [4];
//wire	\eth_udp_inst|ip_send_inst|data_len [5];
//wire	\eth_udp_inst|ip_send_inst|data_len [6];
//wire	\eth_udp_inst|ip_send_inst|data_len [7];
//wire	\eth_udp_inst|ip_send_inst|data_len [8];
//wire	\eth_udp_inst|ip_send_inst|data_len [9];
wire	[3:0] \eth_udp_inst|ip_send_inst|eth_tx_data ;
//wire	\eth_udp_inst|ip_send_inst|eth_tx_data [0];
//wire	\eth_udp_inst|ip_send_inst|eth_tx_data [1];
//wire	\eth_udp_inst|ip_send_inst|eth_tx_data [2];
//wire	\eth_udp_inst|ip_send_inst|eth_tx_data [3];
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~0_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~10_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~11_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~12_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~13_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~14_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~15_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~16_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~17_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~18_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~19_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~1_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~20_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~21_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~22_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~23_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~24_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~25_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~26_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~27_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~28_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~29_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~2_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~30_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~31_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~32_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~33_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~34_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~35_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~36_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~37_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~38_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~39_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~3_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~40_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~41_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~42_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~43_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~44_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~45_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~46_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~47_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~48_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~49_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~4_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~50_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~51_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~52_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~53_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~54_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~55_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~56_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~57_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~58_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~59_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~5_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~60_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~61_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~62_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~63_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~64_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~65_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~66_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~67_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~68_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~69_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~6_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~70_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~71_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~72_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~73_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~74_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~75_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~76_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~77_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~78_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~79_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~7_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~80_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~81_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~82_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~83_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~84_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~85_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~86_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~87_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~88_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~89_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~8_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~90_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~91_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~9_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_en~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~18_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~53_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~21_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~22 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~23_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~24 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~25_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~26 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~27_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~28 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~29_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~30 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~31_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~32 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~33_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~34 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~35_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~36 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~37_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~38 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~39_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~40 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~41_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~42 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~43_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~44 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~45_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~46 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~47_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~48 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~58_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][0]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][10]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][11]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][12]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][13]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][14]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][15]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][1]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][2]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][3]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][4]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][5]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][6]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][7]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][9]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~15_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~17_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~19_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~20_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~49_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~50_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~51_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~52_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~54_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~55_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~56_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~57_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~60_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~61_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~62_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~63_combout ;
wire	\eth_udp_inst|ip_send_inst|packet_head[7][7]~feeder_combout ;
wire	\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ;
wire	\eth_udp_inst|ip_send_inst|read_data_req~0_combout ;
wire	\eth_udp_inst|ip_send_inst|read_data_req~q ;
wire	\eth_udp_inst|ip_send_inst|send_en_r~q ;
wire	\eth_udp_inst|ip_send_inst|send_end~q ;
wire	\eth_udp_inst|ip_send_inst|state.CHECK_SUM~0_combout ;
wire	\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ;
wire	\eth_udp_inst|ip_send_inst|state.CRC~q ;
wire	\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ;
wire	\eth_udp_inst|ip_send_inst|state.IDLE~0_combout ;
wire	\eth_udp_inst|ip_send_inst|state.IDLE~q ;
wire	\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ;
wire	\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ;
wire	\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ;
wire	\eth_udp_inst|ip_send_inst|sw_en~0_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~1_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~2_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~3_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~4_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~5_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~6_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~7_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~q ;
wire	\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X22_Y16_SIG ;
wire	\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ;
wire	\led_r~0_combout ;
wire	\led_r~q ;
wire	[1:0] \mii_to_rmii_inst|eth_tx_data ;
//wire	\mii_to_rmii_inst|eth_tx_data [0];
wire	\mii_to_rmii_inst|eth_tx_data[0]~feeder_combout ;
//wire	\mii_to_rmii_inst|eth_tx_data [1];
wire	[1:0] \mii_to_rmii_inst|eth_tx_data_reg ;
//wire	\mii_to_rmii_inst|eth_tx_data_reg [0];
//wire	\mii_to_rmii_inst|eth_tx_data_reg [1];
wire	\mii_to_rmii_inst|eth_tx_data_reg~0_combout ;
wire	\mii_to_rmii_inst|eth_tx_data_reg~1_combout ;
wire	\mii_to_rmii_inst|eth_tx_dv~feeder_combout ;
wire	\mii_to_rmii_inst|eth_tx_dv~q ;
wire	\mii_to_rmii_inst|rd_flag~0_combout ;
wire	\mii_to_rmii_inst|rd_flag~q ;
wire	[3:0] \mii_to_rmii_inst|tx_data_reg ;
//wire	\mii_to_rmii_inst|tx_data_reg [0];
wire	\mii_to_rmii_inst|tx_data_reg[0]~feeder_combout ;
//wire	\mii_to_rmii_inst|tx_data_reg [1];
wire	\mii_to_rmii_inst|tx_data_reg[1]~feeder_combout ;
//wire	\mii_to_rmii_inst|tx_data_reg [2];
//wire	\mii_to_rmii_inst|tx_data_reg [3];
wire	\mii_to_rmii_inst|tx_data_reg[3]~feeder_combout ;
wire	\mii_to_rmii_inst|tx_dv_reg~feeder_combout ;
wire	\mii_to_rmii_inst|tx_dv_reg~q ;
wire	[5:0] reset_init;
//wire	reset_init[0];
wire	\reset_init[0]~1_combout ;
//wire	reset_init[1];
//wire	reset_init[2];
//wire	reset_init[3];
//wire	reset_init[4];
//wire	reset_init[5];
wire	\reset_init[5]~0_combout ;
wire	\reset_init[5]~clkctrl_outclk ;
wire	\reset_init[5]~clkctrl_outclk__AsyncReset_X17_Y1_INV ;
wire	\rst_n~input_o ;
wire	[24:0] timer;
//wire	timer[0];
wire	\timer[0]~25_combout ;
wire	\timer[0]~26 ;
//wire	timer[10];
wire	\timer[10]~45_combout ;
wire	\timer[10]~46 ;
//wire	timer[11];
wire	\timer[11]~47_combout ;
wire	\timer[11]~48 ;
//wire	timer[12];
wire	\timer[12]~49_combout ;
wire	\timer[12]~50 ;
//wire	timer[13];
wire	\timer[13]~51_combout ;
wire	\timer[13]~52 ;
//wire	timer[14];
wire	\timer[14]~53_combout ;
wire	\timer[14]~54 ;
//wire	timer[15];
wire	\timer[15]~55_combout ;
wire	\timer[15]~56 ;
//wire	timer[16];
wire	\timer[16]~57_combout ;
wire	\timer[16]~58 ;
//wire	timer[17];
wire	\timer[17]~59_combout ;
wire	\timer[17]~60 ;
//wire	timer[18];
wire	\timer[18]~61_combout ;
wire	\timer[18]~62 ;
//wire	timer[19];
wire	\timer[19]~63_combout ;
wire	\timer[19]~64 ;
//wire	timer[1];
wire	\timer[1]~27_combout ;
wire	\timer[1]~28 ;
//wire	timer[20];
wire	\timer[20]~65_combout ;
wire	\timer[20]~66 ;
//wire	timer[21];
wire	\timer[21]~67_combout ;
wire	\timer[21]~68 ;
//wire	timer[22];
wire	\timer[22]~69_combout ;
wire	\timer[22]~70 ;
//wire	timer[23];
wire	\timer[23]~71_combout ;
wire	\timer[23]~72 ;
//wire	timer[24];
wire	\timer[24]~73_combout ;
//wire	timer[2];
wire	\timer[2]~29_combout ;
wire	\timer[2]~30 ;
//wire	timer[3];
wire	\timer[3]~31_combout ;
wire	\timer[3]~32 ;
//wire	timer[4];
wire	\timer[4]~33_combout ;
wire	\timer[4]~34 ;
//wire	timer[5];
wire	\timer[5]~35_combout ;
wire	\timer[5]~36 ;
//wire	timer[6];
wire	\timer[6]~37_combout ;
wire	\timer[6]~38 ;
//wire	timer[7];
wire	\timer[7]~39_combout ;
wire	\timer[7]~40 ;
//wire	timer[8];
wire	\timer[8]~41_combout ;
wire	\timer[8]~42 ;
//wire	timer[9];
wire	\timer[9]~43_combout ;
wire	\timer[9]~44 ;
wire	unknown;

wire vcc;
wire gnd;
assign vcc = 1'b1;
assign gnd = 1'b0;

alta_slice \Add0~8 (
	.A(vcc),
	.B(reset_init[5]),
	.C(vcc),
	.D(vcc),
	.Cin(\Add0~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Add0~8_combout ),
	.Cout(),
	.Q());
defparam \Add0~8 .coord_x = 47;
defparam \Add0~8 .coord_y = 15;
defparam \Add0~8 .coord_z = 12;
defparam \Add0~8 .mask = 16'hC3C3;
defparam \Add0~8 .modeMux = 1'b1;
defparam \Add0~8 .FeedbackMux = 1'b0;
defparam \Add0~8 .ShiftMux = 1'b0;
defparam \Add0~8 .BypassEn = 1'b0;
defparam \Add0~8 .CarryEnb = 1'b1;

alta_slice \Equal0~0 (
	.A(timer[1]),
	.B(timer[3]),
	.C(timer[2]),
	.D(timer[0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~0_combout ),
	.Cout(),
	.Q());
defparam \Equal0~0 .coord_x = 2;
defparam \Equal0~0 .coord_y = 10;
defparam \Equal0~0 .coord_z = 0;
defparam \Equal0~0 .mask = 16'h0001;
defparam \Equal0~0 .modeMux = 1'b0;
defparam \Equal0~0 .FeedbackMux = 1'b0;
defparam \Equal0~0 .ShiftMux = 1'b0;
defparam \Equal0~0 .BypassEn = 1'b0;
defparam \Equal0~0 .CarryEnb = 1'b1;

alta_slice \Equal0~1 (
	.A(timer[7]),
	.B(timer[5]),
	.C(timer[6]),
	.D(timer[4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~1_combout ),
	.Cout(),
	.Q());
defparam \Equal0~1 .coord_x = 2;
defparam \Equal0~1 .coord_y = 10;
defparam \Equal0~1 .coord_z = 1;
defparam \Equal0~1 .mask = 16'h0001;
defparam \Equal0~1 .modeMux = 1'b0;
defparam \Equal0~1 .FeedbackMux = 1'b0;
defparam \Equal0~1 .ShiftMux = 1'b0;
defparam \Equal0~1 .BypassEn = 1'b0;
defparam \Equal0~1 .CarryEnb = 1'b1;

alta_slice \Equal0~2 (
	.A(timer[11]),
	.B(timer[10]),
	.C(timer[8]),
	.D(timer[9]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~2_combout ),
	.Cout(),
	.Q());
defparam \Equal0~2 .coord_x = 2;
defparam \Equal0~2 .coord_y = 10;
defparam \Equal0~2 .coord_z = 2;
defparam \Equal0~2 .mask = 16'h0001;
defparam \Equal0~2 .modeMux = 1'b0;
defparam \Equal0~2 .FeedbackMux = 1'b0;
defparam \Equal0~2 .ShiftMux = 1'b0;
defparam \Equal0~2 .BypassEn = 1'b0;
defparam \Equal0~2 .CarryEnb = 1'b1;

alta_slice \Equal0~3 (
	.A(timer[13]),
	.B(timer[14]),
	.C(timer[15]),
	.D(timer[12]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~3_combout ),
	.Cout(),
	.Q());
defparam \Equal0~3 .coord_x = 2;
defparam \Equal0~3 .coord_y = 9;
defparam \Equal0~3 .coord_z = 13;
defparam \Equal0~3 .mask = 16'h0001;
defparam \Equal0~3 .modeMux = 1'b0;
defparam \Equal0~3 .FeedbackMux = 1'b0;
defparam \Equal0~3 .ShiftMux = 1'b0;
defparam \Equal0~3 .BypassEn = 1'b0;
defparam \Equal0~3 .CarryEnb = 1'b1;

alta_slice \Equal0~4 (
	.A(\Equal0~0_combout ),
	.B(\Equal0~2_combout ),
	.C(\Equal0~1_combout ),
	.D(\Equal0~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~4_combout ),
	.Cout(),
	.Q());
defparam \Equal0~4 .coord_x = 2;
defparam \Equal0~4 .coord_y = 10;
defparam \Equal0~4 .coord_z = 3;
defparam \Equal0~4 .mask = 16'h8000;
defparam \Equal0~4 .modeMux = 1'b0;
defparam \Equal0~4 .FeedbackMux = 1'b0;
defparam \Equal0~4 .ShiftMux = 1'b0;
defparam \Equal0~4 .BypassEn = 1'b0;
defparam \Equal0~4 .CarryEnb = 1'b1;

alta_slice \Equal0~5 (
	.A(timer[17]),
	.B(timer[19]),
	.C(timer[16]),
	.D(timer[18]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~5_combout ),
	.Cout(),
	.Q());
defparam \Equal0~5 .coord_x = 2;
defparam \Equal0~5 .coord_y = 9;
defparam \Equal0~5 .coord_z = 14;
defparam \Equal0~5 .mask = 16'h0001;
defparam \Equal0~5 .modeMux = 1'b0;
defparam \Equal0~5 .FeedbackMux = 1'b0;
defparam \Equal0~5 .ShiftMux = 1'b0;
defparam \Equal0~5 .BypassEn = 1'b0;
defparam \Equal0~5 .CarryEnb = 1'b1;

alta_slice \Equal0~6 (
	.A(timer[23]),
	.B(timer[20]),
	.C(timer[21]),
	.D(timer[22]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~6_combout ),
	.Cout(),
	.Q());
defparam \Equal0~6 .coord_x = 2;
defparam \Equal0~6 .coord_y = 9;
defparam \Equal0~6 .coord_z = 15;
defparam \Equal0~6 .mask = 16'h0001;
defparam \Equal0~6 .modeMux = 1'b0;
defparam \Equal0~6 .FeedbackMux = 1'b0;
defparam \Equal0~6 .ShiftMux = 1'b0;
defparam \Equal0~6 .BypassEn = 1'b0;
defparam \Equal0~6 .CarryEnb = 1'b1;

alta_slice \Equal0~7 (
	.A(vcc),
	.B(vcc),
	.C(\Equal0~6_combout ),
	.D(timer[24]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~7_combout ),
	.Cout(),
	.Q());
defparam \Equal0~7 .coord_x = 1;
defparam \Equal0~7 .coord_y = 9;
defparam \Equal0~7 .coord_z = 13;
defparam \Equal0~7 .mask = 16'h00F0;
defparam \Equal0~7 .modeMux = 1'b0;
defparam \Equal0~7 .FeedbackMux = 1'b0;
defparam \Equal0~7 .ShiftMux = 1'b0;
defparam \Equal0~7 .BypassEn = 1'b0;
defparam \Equal0~7 .CarryEnb = 1'b1;

alta_slice \alt_pll_inst|altpll_component|auto_generated|locked (
	.A(\alt_pll_inst|altpll_component|auto_generated|pll_lock_sync~q ),
	.B(vcc),
	.C(vcc),
	.D(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.Cout(),
	.Q());
defparam \alt_pll_inst|altpll_component|auto_generated|locked .coord_x = 1;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .coord_y = 1;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .coord_z = 9;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .mask = 16'h55FF;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .modeMux = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .FeedbackMux = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .ShiftMux = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .BypassEn = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .CarryEnb = 1'b1;

alta_io_gclk \alt_pll_inst|altpll_component|auto_generated|locked~clkctrl (
	.inclk(\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.outclk(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ));
defparam \alt_pll_inst|altpll_component|auto_generated|locked~clkctrl .coord_x = 49;
defparam \alt_pll_inst|altpll_component|auto_generated|locked~clkctrl .coord_y = 15;
defparam \alt_pll_inst|altpll_component|auto_generated|locked~clkctrl .coord_z = 2;

alta_pllve \alt_pll_inst|altpll_component|auto_generated|pll1 (
	.clkin(\clk~input_o ),
	.clkfb(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_fbout ),
	.pfden(vcc),
	.resetn(\reset_init[5]~clkctrl_outclk ),
	.phasecounterselect({gnd, gnd, gnd}),
	.phaseupdown(gnd),
	.phasestep(gnd),
	.scanclk(gnd),
	.scanclkena(vcc),
	.scandata(gnd),
	.configupdate(gnd),
	.scandataout(),
	.scandone(),
	.phasedone(),
	.clkout0(\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [0]),
	.clkout1(\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [1]),
	.clkout2(\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [2]),
	.clkout3(\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [3]),
	.clkout4(\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [4]),
	.clkfbout(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_fbout ),
	.lock(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked ));
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .coord_x = 0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .coord_y = 1;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .coord_z = 0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKIN_HIGH = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKIN_LOW = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKIN_TRIM = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKIN_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKFB_HIGH = 8'b00010001;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKFB_LOW = 8'b00010010;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKFB_TRIM = 1'b1;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKFB_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKDIV0_EN = 1'b1;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKDIV1_EN = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKDIV2_EN = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKDIV3_EN = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKDIV4_EN = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT0_HIGH = 8'b00010001;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT0_LOW = 8'b00010010;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT0_TRIM = 1'b1;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT0_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_HIGH = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_LOW = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_TRIM = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_HIGH = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_LOW = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_TRIM = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_HIGH = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_LOW = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_TRIM = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_HIGH = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_LOW = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_TRIM = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT0_DEL = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_DEL = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_DEL = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_DEL = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_DEL = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT0_PHASE = 3'b000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_PHASE = 3'b000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_PHASE = 3'b000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_PHASE = 3'b000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_PHASE = 3'b000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKFB_DEL = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKFB_PHASE = 3'b000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .FEEDBACK_MODE = 3'b100;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .FBDELAY_VAL = 3'b100;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .PLLOUTP_EN = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .PLLOUTN_EN = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_CASCADE = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_CASCADE = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_CASCADE = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_CASCADE = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .VCO_POST_DIV = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .REG_CTRL = 2'b10;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CP = 3'b100;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .RREF = 2'b01;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .RVI = 2'b01;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .IVCO = 3'b010;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .PLL_EN_FLAG = 1'b1;

alta_slice \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\alt_pll_inst|altpll_component|auto_generated|pll_lock_sync~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked_X17_Y1_SIG_VCC ),
	.AsyncReset(\reset_init[5]~clkctrl_outclk__AsyncReset_X17_Y1_INV ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\alt_pll_inst|altpll_component|auto_generated|pll_lock_sync~feeder_combout ),
	.Cout(),
	.Q(\alt_pll_inst|altpll_component|auto_generated|pll_lock_sync~q ));
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .coord_x = 1;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .coord_y = 1;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .coord_z = 3;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .mask = 16'hFFFF;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .modeMux = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .FeedbackMux = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .ShiftMux = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .BypassEn = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .CarryEnb = 1'b1;

alta_io_gclk \alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl (
	.inclk(\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [0]),
	.outclk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ));
defparam \alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl .coord_x = 0;
defparam \alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl .coord_y = 12;
defparam \alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl .coord_z = 3;

alta_asyncctrl asyncreset_ctrl_X11_Y15_N0(
	.Din(),
	.Dout(AsyncReset_X11_Y15_GND));
defparam asyncreset_ctrl_X11_Y15_N0.coord_x = 1;
defparam asyncreset_ctrl_X11_Y15_N0.coord_y = 9;
defparam asyncreset_ctrl_X11_Y15_N0.coord_z = 0;
defparam asyncreset_ctrl_X11_Y15_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X12_Y12_N0(
	.Din(),
	.Dout(AsyncReset_X12_Y12_GND));
defparam asyncreset_ctrl_X12_Y12_N0.coord_x = 47;
defparam asyncreset_ctrl_X12_Y12_N0.coord_y = 15;
defparam asyncreset_ctrl_X12_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X12_Y12_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X12_Y13_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ));
defparam asyncreset_ctrl_X12_Y13_N0.coord_x = 16;
defparam asyncreset_ctrl_X12_Y13_N0.coord_y = 13;
defparam asyncreset_ctrl_X12_Y13_N0.coord_z = 0;
defparam asyncreset_ctrl_X12_Y13_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X12_Y14_N0(
	.Din(),
	.Dout(AsyncReset_X12_Y14_GND));
defparam asyncreset_ctrl_X12_Y14_N0.coord_x = 2;
defparam asyncreset_ctrl_X12_Y14_N0.coord_y = 9;
defparam asyncreset_ctrl_X12_Y14_N0.coord_z = 0;
defparam asyncreset_ctrl_X12_Y14_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X12_Y15_N0(
	.Din(),
	.Dout(AsyncReset_X12_Y15_GND));
defparam asyncreset_ctrl_X12_Y15_N0.coord_x = 2;
defparam asyncreset_ctrl_X12_Y15_N0.coord_y = 10;
defparam asyncreset_ctrl_X12_Y15_N0.coord_z = 0;
defparam asyncreset_ctrl_X12_Y15_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X13_Y12_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ));
defparam asyncreset_ctrl_X13_Y12_N0.coord_x = 15;
defparam asyncreset_ctrl_X13_Y12_N0.coord_y = 16;
defparam asyncreset_ctrl_X13_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X13_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X13_Y13_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y13_SIG ));
defparam asyncreset_ctrl_X13_Y13_N0.coord_x = 15;
defparam asyncreset_ctrl_X13_Y13_N0.coord_y = 13;
defparam asyncreset_ctrl_X13_Y13_N0.coord_z = 0;
defparam asyncreset_ctrl_X13_Y13_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X14_Y12_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y12_SIG ));
defparam asyncreset_ctrl_X14_Y12_N0.coord_x = 17;
defparam asyncreset_ctrl_X14_Y12_N0.coord_y = 16;
defparam asyncreset_ctrl_X14_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X14_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X14_Y13_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ));
defparam asyncreset_ctrl_X14_Y13_N0.coord_x = 17;
defparam asyncreset_ctrl_X14_Y13_N0.coord_y = 13;
defparam asyncreset_ctrl_X14_Y13_N0.coord_z = 0;
defparam asyncreset_ctrl_X14_Y13_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X14_Y17_N1(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X14_Y17_SIG ));
defparam asyncreset_ctrl_X14_Y17_N1.coord_x = 10;
defparam asyncreset_ctrl_X14_Y17_N1.coord_y = 15;
defparam asyncreset_ctrl_X14_Y17_N1.coord_z = 1;
defparam asyncreset_ctrl_X14_Y17_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X16_Y11_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ));
defparam asyncreset_ctrl_X16_Y11_N0.coord_x = 17;
defparam asyncreset_ctrl_X16_Y11_N0.coord_y = 15;
defparam asyncreset_ctrl_X16_Y11_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y11_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X16_Y12_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ));
defparam asyncreset_ctrl_X16_Y12_N0.coord_x = 16;
defparam asyncreset_ctrl_X16_Y12_N0.coord_y = 16;
defparam asyncreset_ctrl_X16_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X16_Y13_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ));
defparam asyncreset_ctrl_X16_Y13_N0.coord_x = 17;
defparam asyncreset_ctrl_X16_Y13_N0.coord_y = 14;
defparam asyncreset_ctrl_X16_Y13_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y13_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X16_Y16_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y16_SIG ));
defparam asyncreset_ctrl_X16_Y16_N0.coord_x = 11;
defparam asyncreset_ctrl_X16_Y16_N0.coord_y = 15;
defparam asyncreset_ctrl_X16_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y16_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X16_Y17_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y17_SIG ));
defparam asyncreset_ctrl_X16_Y17_N0.coord_x = 10;
defparam asyncreset_ctrl_X16_Y17_N0.coord_y = 13;
defparam asyncreset_ctrl_X16_Y17_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y17_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X16_Y18_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y18_SIG ));
defparam asyncreset_ctrl_X16_Y18_N0.coord_x = 11;
defparam asyncreset_ctrl_X16_Y18_N0.coord_y = 14;
defparam asyncreset_ctrl_X16_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y18_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X17_Y12_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y12_SIG ));
defparam asyncreset_ctrl_X17_Y12_N0.coord_x = 15;
defparam asyncreset_ctrl_X17_Y12_N0.coord_y = 15;
defparam asyncreset_ctrl_X17_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X17_Y13_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ));
defparam asyncreset_ctrl_X17_Y13_N0.coord_x = 16;
defparam asyncreset_ctrl_X17_Y13_N0.coord_y = 15;
defparam asyncreset_ctrl_X17_Y13_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y13_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X17_Y14_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y14_SIG ));
defparam asyncreset_ctrl_X17_Y14_N0.coord_x = 16;
defparam asyncreset_ctrl_X17_Y14_N0.coord_y = 14;
defparam asyncreset_ctrl_X17_Y14_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y14_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X17_Y17_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y17_SIG ));
defparam asyncreset_ctrl_X17_Y17_N0.coord_x = 11;
defparam asyncreset_ctrl_X17_Y17_N0.coord_y = 13;
defparam asyncreset_ctrl_X17_Y17_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y17_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X17_Y1_N0(
	.Din(\reset_init[5]~clkctrl_outclk ),
	.Dout(\reset_init[5]~clkctrl_outclk__AsyncReset_X17_Y1_INV ));
defparam asyncreset_ctrl_X17_Y1_N0.coord_x = 1;
defparam asyncreset_ctrl_X17_Y1_N0.coord_y = 1;
defparam asyncreset_ctrl_X17_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y1_N0.AsyncCtrlMux = 2'b11;

alta_asyncctrl asyncreset_ctrl_X18_Y17_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y17_SIG ));
defparam asyncreset_ctrl_X18_Y17_N0.coord_x = 13;
defparam asyncreset_ctrl_X18_Y17_N0.coord_y = 13;
defparam asyncreset_ctrl_X18_Y17_N0.coord_z = 0;
defparam asyncreset_ctrl_X18_Y17_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X19_Y12_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X19_Y12_SIG ));
defparam asyncreset_ctrl_X19_Y12_N0.coord_x = 19;
defparam asyncreset_ctrl_X19_Y12_N0.coord_y = 16;
defparam asyncreset_ctrl_X19_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X19_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X1_Y17_N1(
	.Din(),
	.Dout(AsyncReset_X1_Y17_GND));
defparam asyncreset_ctrl_X1_Y17_N1.coord_x = 11;
defparam asyncreset_ctrl_X1_Y17_N1.coord_y = 16;
defparam asyncreset_ctrl_X1_Y17_N1.coord_z = 1;
defparam asyncreset_ctrl_X1_Y17_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X1_Y7_N0(
	.Din(),
	.Dout(AsyncReset_X1_Y7_GND));
defparam asyncreset_ctrl_X1_Y7_N0.coord_x = 8;
defparam asyncreset_ctrl_X1_Y7_N0.coord_y = 12;
defparam asyncreset_ctrl_X1_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X1_Y7_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X21_Y18_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ));
defparam asyncreset_ctrl_X21_Y18_N0.coord_x = 20;
defparam asyncreset_ctrl_X21_Y18_N0.coord_y = 16;
defparam asyncreset_ctrl_X21_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X21_Y18_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X21_Y19_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y19_SIG ));
defparam asyncreset_ctrl_X21_Y19_N0.coord_x = 20;
defparam asyncreset_ctrl_X21_Y19_N0.coord_y = 17;
defparam asyncreset_ctrl_X21_Y19_N0.coord_z = 0;
defparam asyncreset_ctrl_X21_Y19_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X22_Y16_N1(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y16_SIG ));
defparam asyncreset_ctrl_X22_Y16_N1.coord_x = 22;
defparam asyncreset_ctrl_X22_Y16_N1.coord_y = 16;
defparam asyncreset_ctrl_X22_Y16_N1.coord_z = 1;
defparam asyncreset_ctrl_X22_Y16_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X22_Y19_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ));
defparam asyncreset_ctrl_X22_Y19_N0.coord_x = 19;
defparam asyncreset_ctrl_X22_Y19_N0.coord_y = 17;
defparam asyncreset_ctrl_X22_Y19_N0.coord_z = 0;
defparam asyncreset_ctrl_X22_Y19_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X22_Y8_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y8_SIG ));
defparam asyncreset_ctrl_X22_Y8_N0.coord_x = 10;
defparam asyncreset_ctrl_X22_Y8_N0.coord_y = 17;
defparam asyncreset_ctrl_X22_Y8_N0.coord_z = 0;
defparam asyncreset_ctrl_X22_Y8_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X23_Y15_N1(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ));
defparam asyncreset_ctrl_X23_Y15_N1.coord_x = 22;
defparam asyncreset_ctrl_X23_Y15_N1.coord_y = 18;
defparam asyncreset_ctrl_X23_Y15_N1.coord_z = 1;
defparam asyncreset_ctrl_X23_Y15_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X23_Y16_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ));
defparam asyncreset_ctrl_X23_Y16_N0.coord_x = 21;
defparam asyncreset_ctrl_X23_Y16_N0.coord_y = 13;
defparam asyncreset_ctrl_X23_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X23_Y16_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X23_Y18_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y18_SIG ));
defparam asyncreset_ctrl_X23_Y18_N0.coord_x = 21;
defparam asyncreset_ctrl_X23_Y18_N0.coord_y = 16;
defparam asyncreset_ctrl_X23_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X23_Y18_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X23_Y19_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y19_SIG ));
defparam asyncreset_ctrl_X23_Y19_N0.coord_x = 21;
defparam asyncreset_ctrl_X23_Y19_N0.coord_y = 17;
defparam asyncreset_ctrl_X23_Y19_N0.coord_z = 0;
defparam asyncreset_ctrl_X23_Y19_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X23_Y8_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ));
defparam asyncreset_ctrl_X23_Y8_N0.coord_x = 11;
defparam asyncreset_ctrl_X23_Y8_N0.coord_y = 17;
defparam asyncreset_ctrl_X23_Y8_N0.coord_z = 0;
defparam asyncreset_ctrl_X23_Y8_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X24_Y15_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ));
defparam asyncreset_ctrl_X24_Y15_N0.coord_x = 20;
defparam asyncreset_ctrl_X24_Y15_N0.coord_y = 15;
defparam asyncreset_ctrl_X24_Y15_N0.coord_z = 0;
defparam asyncreset_ctrl_X24_Y15_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X24_Y15_N1(
	.Din(),
	.Dout(AsyncReset_X24_Y15_GND));
defparam asyncreset_ctrl_X24_Y15_N1.coord_x = 20;
defparam asyncreset_ctrl_X24_Y15_N1.coord_y = 15;
defparam asyncreset_ctrl_X24_Y15_N1.coord_z = 1;
defparam asyncreset_ctrl_X24_Y15_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X24_Y16_N1(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ));
defparam asyncreset_ctrl_X24_Y16_N1.coord_x = 22;
defparam asyncreset_ctrl_X24_Y16_N1.coord_y = 14;
defparam asyncreset_ctrl_X24_Y16_N1.coord_z = 1;
defparam asyncreset_ctrl_X24_Y16_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X25_Y16_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y16_SIG ));
defparam asyncreset_ctrl_X25_Y16_N0.coord_x = 21;
defparam asyncreset_ctrl_X25_Y16_N0.coord_y = 14;
defparam asyncreset_ctrl_X25_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X25_Y16_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X25_Y17_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ));
defparam asyncreset_ctrl_X25_Y17_N0.coord_x = 19;
defparam asyncreset_ctrl_X25_Y17_N0.coord_y = 11;
defparam asyncreset_ctrl_X25_Y17_N0.coord_z = 0;
defparam asyncreset_ctrl_X25_Y17_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X28_Y14_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y14_SIG ));
defparam asyncreset_ctrl_X28_Y14_N0.coord_x = 21;
defparam asyncreset_ctrl_X28_Y14_N0.coord_y = 9;
defparam asyncreset_ctrl_X28_Y14_N0.coord_z = 0;
defparam asyncreset_ctrl_X28_Y14_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X28_Y14_N1(
	.Din(),
	.Dout(AsyncReset_X28_Y14_GND));
defparam asyncreset_ctrl_X28_Y14_N1.coord_x = 21;
defparam asyncreset_ctrl_X28_Y14_N1.coord_y = 9;
defparam asyncreset_ctrl_X28_Y14_N1.coord_z = 1;
defparam asyncreset_ctrl_X28_Y14_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X28_Y15_N0(
	.Din(),
	.Dout(AsyncReset_X28_Y15_GND));
defparam asyncreset_ctrl_X28_Y15_N0.coord_x = 21;
defparam asyncreset_ctrl_X28_Y15_N0.coord_y = 10;
defparam asyncreset_ctrl_X28_Y15_N0.coord_z = 0;
defparam asyncreset_ctrl_X28_Y15_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X28_Y15_N1(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y15_SIG ));
defparam asyncreset_ctrl_X28_Y15_N1.coord_x = 21;
defparam asyncreset_ctrl_X28_Y15_N1.coord_y = 10;
defparam asyncreset_ctrl_X28_Y15_N1.coord_z = 1;
defparam asyncreset_ctrl_X28_Y15_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X28_Y18_N0(
	.Din(),
	.Dout(AsyncReset_X28_Y18_GND));
defparam asyncreset_ctrl_X28_Y18_N0.coord_x = 20;
defparam asyncreset_ctrl_X28_Y18_N0.coord_y = 10;
defparam asyncreset_ctrl_X28_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X28_Y18_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X2_Y7_N0(
	.Din(),
	.Dout(AsyncReset_X2_Y7_GND));
defparam asyncreset_ctrl_X2_Y7_N0.coord_x = 9;
defparam asyncreset_ctrl_X2_Y7_N0.coord_y = 12;
defparam asyncreset_ctrl_X2_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X2_Y7_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X33_Y15_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y15_SIG ));
defparam asyncreset_ctrl_X33_Y15_N0.coord_x = 46;
defparam asyncreset_ctrl_X33_Y15_N0.coord_y = 15;
defparam asyncreset_ctrl_X33_Y15_N0.coord_z = 0;
defparam asyncreset_ctrl_X33_Y15_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X3_Y7_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X3_Y7_SIG ));
defparam asyncreset_ctrl_X3_Y7_N0.coord_x = 14;
defparam asyncreset_ctrl_X3_Y7_N0.coord_y = 16;
defparam asyncreset_ctrl_X3_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X3_Y7_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X4_Y7_N0(
	.Din(),
	.Dout(AsyncReset_X4_Y7_GND));
defparam asyncreset_ctrl_X4_Y7_N0.coord_x = 17;
defparam asyncreset_ctrl_X4_Y7_N0.coord_y = 12;
defparam asyncreset_ctrl_X4_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X4_Y7_N0.AsyncCtrlMux = 2'b00;

alta_dio \cam_data[0]~input (
	.padio(cam_data[0]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[0]~input_o ),
	.regout());
defparam \cam_data[0]~input .coord_x = 11;
defparam \cam_data[0]~input .coord_y = 0;
defparam \cam_data[0]~input .coord_z = 1;
defparam \cam_data[0]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[0]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[0]~input .IN_POWERUP = 1'b0;
defparam \cam_data[0]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[0]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[0]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[0]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[0]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[0]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[0]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[0]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[0]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[0]~input .OUT_DDIO = 1'b0;
defparam \cam_data[0]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[0]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[0]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[0]~input .OE_POWERUP = 1'b0;
defparam \cam_data[0]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[0]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[0]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[0]~input .OE_DDIO = 1'b0;
defparam \cam_data[0]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[0]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[0]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[0]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[0]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[0]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[0]~input .CFG_KEEP = 2'b00;
defparam \cam_data[0]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[0]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[0]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[0]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[0]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[0]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[0]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[0]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[0]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[0]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[0]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[0]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[0]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[0]~input .OUT_DELAY = 1'b0;
defparam \cam_data[0]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[0]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[1]~input (
	.padio(cam_data[1]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[1]~input_o ),
	.regout());
defparam \cam_data[1]~input .coord_x = 6;
defparam \cam_data[1]~input .coord_y = 0;
defparam \cam_data[1]~input .coord_z = 0;
defparam \cam_data[1]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[1]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[1]~input .IN_POWERUP = 1'b0;
defparam \cam_data[1]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[1]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[1]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[1]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[1]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[1]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[1]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[1]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[1]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[1]~input .OUT_DDIO = 1'b0;
defparam \cam_data[1]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[1]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[1]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[1]~input .OE_POWERUP = 1'b0;
defparam \cam_data[1]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[1]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[1]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[1]~input .OE_DDIO = 1'b0;
defparam \cam_data[1]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[1]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[1]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[1]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[1]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[1]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[1]~input .CFG_KEEP = 2'b00;
defparam \cam_data[1]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[1]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[1]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[1]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[1]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[1]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[1]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[1]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[1]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[1]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[1]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[1]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[1]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[1]~input .OUT_DELAY = 1'b0;
defparam \cam_data[1]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[1]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[2]~input (
	.padio(cam_data[2]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[2]~input_o ),
	.regout());
defparam \cam_data[2]~input .coord_x = 6;
defparam \cam_data[2]~input .coord_y = 0;
defparam \cam_data[2]~input .coord_z = 1;
defparam \cam_data[2]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[2]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[2]~input .IN_POWERUP = 1'b0;
defparam \cam_data[2]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[2]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[2]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[2]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[2]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[2]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[2]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[2]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[2]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[2]~input .OUT_DDIO = 1'b0;
defparam \cam_data[2]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[2]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[2]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[2]~input .OE_POWERUP = 1'b0;
defparam \cam_data[2]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[2]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[2]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[2]~input .OE_DDIO = 1'b0;
defparam \cam_data[2]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[2]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[2]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[2]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[2]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[2]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[2]~input .CFG_KEEP = 2'b00;
defparam \cam_data[2]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[2]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[2]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[2]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[2]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[2]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[2]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[2]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[2]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[2]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[2]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[2]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[2]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[2]~input .OUT_DELAY = 1'b0;
defparam \cam_data[2]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[2]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[3]~input (
	.padio(cam_data[3]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[3]~input_o ),
	.regout());
defparam \cam_data[3]~input .coord_x = 5;
defparam \cam_data[3]~input .coord_y = 0;
defparam \cam_data[3]~input .coord_z = 2;
defparam \cam_data[3]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[3]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[3]~input .IN_POWERUP = 1'b0;
defparam \cam_data[3]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[3]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[3]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[3]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[3]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[3]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[3]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[3]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[3]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[3]~input .OUT_DDIO = 1'b0;
defparam \cam_data[3]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[3]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[3]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[3]~input .OE_POWERUP = 1'b0;
defparam \cam_data[3]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[3]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[3]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[3]~input .OE_DDIO = 1'b0;
defparam \cam_data[3]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[3]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[3]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[3]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[3]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[3]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[3]~input .CFG_KEEP = 2'b00;
defparam \cam_data[3]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[3]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[3]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[3]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[3]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[3]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[3]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[3]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[3]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[3]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[3]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[3]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[3]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[3]~input .OUT_DELAY = 1'b0;
defparam \cam_data[3]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[3]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[4]~input (
	.padio(cam_data[4]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[4]~input_o ),
	.regout());
defparam \cam_data[4]~input .coord_x = 3;
defparam \cam_data[4]~input .coord_y = 0;
defparam \cam_data[4]~input .coord_z = 0;
defparam \cam_data[4]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[4]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[4]~input .IN_POWERUP = 1'b0;
defparam \cam_data[4]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[4]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[4]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[4]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[4]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[4]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[4]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[4]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[4]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[4]~input .OUT_DDIO = 1'b0;
defparam \cam_data[4]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[4]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[4]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[4]~input .OE_POWERUP = 1'b0;
defparam \cam_data[4]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[4]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[4]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[4]~input .OE_DDIO = 1'b0;
defparam \cam_data[4]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[4]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[4]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[4]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[4]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[4]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[4]~input .CFG_KEEP = 2'b00;
defparam \cam_data[4]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[4]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[4]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[4]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[4]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[4]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[4]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[4]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[4]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[4]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[4]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[4]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[4]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[4]~input .OUT_DELAY = 1'b0;
defparam \cam_data[4]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[4]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[5]~input (
	.padio(cam_data[5]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[5]~input_o ),
	.regout());
defparam \cam_data[5]~input .coord_x = 3;
defparam \cam_data[5]~input .coord_y = 0;
defparam \cam_data[5]~input .coord_z = 1;
defparam \cam_data[5]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[5]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[5]~input .IN_POWERUP = 1'b0;
defparam \cam_data[5]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[5]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[5]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[5]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[5]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[5]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[5]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[5]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[5]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[5]~input .OUT_DDIO = 1'b0;
defparam \cam_data[5]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[5]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[5]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[5]~input .OE_POWERUP = 1'b0;
defparam \cam_data[5]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[5]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[5]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[5]~input .OE_DDIO = 1'b0;
defparam \cam_data[5]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[5]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[5]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[5]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[5]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[5]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[5]~input .CFG_KEEP = 2'b00;
defparam \cam_data[5]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[5]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[5]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[5]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[5]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[5]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[5]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[5]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[5]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[5]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[5]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[5]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[5]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[5]~input .OUT_DELAY = 1'b0;
defparam \cam_data[5]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[5]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[6]~input (
	.padio(cam_data[6]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[6]~input_o ),
	.regout());
defparam \cam_data[6]~input .coord_x = 0;
defparam \cam_data[6]~input .coord_y = 4;
defparam \cam_data[6]~input .coord_z = 2;
defparam \cam_data[6]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[6]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[6]~input .IN_POWERUP = 1'b0;
defparam \cam_data[6]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[6]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[6]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[6]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[6]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[6]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[6]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[6]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[6]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[6]~input .OUT_DDIO = 1'b0;
defparam \cam_data[6]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[6]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[6]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[6]~input .OE_POWERUP = 1'b0;
defparam \cam_data[6]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[6]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[6]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[6]~input .OE_DDIO = 1'b0;
defparam \cam_data[6]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[6]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[6]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[6]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[6]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[6]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[6]~input .CFG_KEEP = 2'b00;
defparam \cam_data[6]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[6]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[6]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[6]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[6]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[6]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[6]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[6]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[6]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[6]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[6]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[6]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[6]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[6]~input .OUT_DELAY = 1'b0;
defparam \cam_data[6]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[6]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[7]~input (
	.padio(cam_data[7]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[7]~input_o ),
	.regout());
defparam \cam_data[7]~input .coord_x = 0;
defparam \cam_data[7]~input .coord_y = 4;
defparam \cam_data[7]~input .coord_z = 3;
defparam \cam_data[7]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[7]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[7]~input .IN_POWERUP = 1'b0;
defparam \cam_data[7]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[7]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[7]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[7]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[7]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[7]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[7]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[7]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[7]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[7]~input .OUT_DDIO = 1'b0;
defparam \cam_data[7]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[7]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[7]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[7]~input .OE_POWERUP = 1'b0;
defparam \cam_data[7]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[7]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[7]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[7]~input .OE_DDIO = 1'b0;
defparam \cam_data[7]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[7]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[7]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[7]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[7]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[7]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[7]~input .CFG_KEEP = 2'b00;
defparam \cam_data[7]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[7]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[7]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[7]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[7]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[7]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[7]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[7]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[7]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[7]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[7]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[7]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[7]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[7]~input .OUT_DELAY = 1'b0;
defparam \cam_data[7]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[7]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_hsync~input (
	.padio(cam_hsync),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_hsync~input_o ),
	.regout());
defparam \cam_hsync~input .coord_x = 0;
defparam \cam_hsync~input .coord_y = 8;
defparam \cam_hsync~input .coord_z = 2;
defparam \cam_hsync~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_hsync~input .IN_SYNC_MODE = 1'b0;
defparam \cam_hsync~input .IN_POWERUP = 1'b0;
defparam \cam_hsync~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_hsync~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_hsync~input .OUT_REG_MODE = 1'b0;
defparam \cam_hsync~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_hsync~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_hsync~input .OUT_POWERUP = 1'b0;
defparam \cam_hsync~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_hsync~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_hsync~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_hsync~input .OUT_DDIO = 1'b0;
defparam \cam_hsync~input .OE_REG_MODE = 1'b0;
defparam \cam_hsync~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_hsync~input .OE_SYNC_MODE = 1'b0;
defparam \cam_hsync~input .OE_POWERUP = 1'b0;
defparam \cam_hsync~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_hsync~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_hsync~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_hsync~input .OE_DDIO = 1'b0;
defparam \cam_hsync~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_hsync~input .CFG_PULL_UP = 1'b0;
defparam \cam_hsync~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_hsync~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_hsync~input .CFG_PDRV = 7'b0011010;
defparam \cam_hsync~input .CFG_NDRV = 7'b0011000;
defparam \cam_hsync~input .CFG_KEEP = 2'b00;
defparam \cam_hsync~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_hsync~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_hsync~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_hsync~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_hsync~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_hsync~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_hsync~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_hsync~input .CFG_OSCDIV = 2'b00;
defparam \cam_hsync~input .CFG_ROCTUSR = 1'b0;
defparam \cam_hsync~input .CFG_SEL_CUA = 1'b0;
defparam \cam_hsync~input .CFG_ROCT_EN = 1'b0;
defparam \cam_hsync~input .INPUT_ONLY = 1'b0;
defparam \cam_hsync~input .DPCLK_DELAY = 4'b0000;
defparam \cam_hsync~input .OUT_DELAY = 1'b0;
defparam \cam_hsync~input .IN_DATA_DELAY = 3'b000;
defparam \cam_hsync~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_pclk~input (
	.padio(cam_pclk),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_pclk~input_o ),
	.regout());
defparam \cam_pclk~input .coord_x = 0;
defparam \cam_pclk~input .coord_y = 8;
defparam \cam_pclk~input .coord_z = 1;
defparam \cam_pclk~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_pclk~input .IN_SYNC_MODE = 1'b0;
defparam \cam_pclk~input .IN_POWERUP = 1'b0;
defparam \cam_pclk~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_pclk~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_pclk~input .OUT_REG_MODE = 1'b0;
defparam \cam_pclk~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_pclk~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_pclk~input .OUT_POWERUP = 1'b0;
defparam \cam_pclk~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_pclk~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_pclk~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_pclk~input .OUT_DDIO = 1'b0;
defparam \cam_pclk~input .OE_REG_MODE = 1'b0;
defparam \cam_pclk~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_pclk~input .OE_SYNC_MODE = 1'b0;
defparam \cam_pclk~input .OE_POWERUP = 1'b0;
defparam \cam_pclk~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_pclk~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_pclk~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_pclk~input .OE_DDIO = 1'b0;
defparam \cam_pclk~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_pclk~input .CFG_PULL_UP = 1'b0;
defparam \cam_pclk~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_pclk~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_pclk~input .CFG_PDRV = 7'b0011010;
defparam \cam_pclk~input .CFG_NDRV = 7'b0011000;
defparam \cam_pclk~input .CFG_KEEP = 2'b00;
defparam \cam_pclk~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_pclk~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_pclk~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_pclk~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_pclk~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_pclk~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_pclk~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_pclk~input .CFG_OSCDIV = 2'b00;
defparam \cam_pclk~input .CFG_ROCTUSR = 1'b0;
defparam \cam_pclk~input .CFG_SEL_CUA = 1'b0;
defparam \cam_pclk~input .CFG_ROCT_EN = 1'b0;
defparam \cam_pclk~input .INPUT_ONLY = 1'b0;
defparam \cam_pclk~input .DPCLK_DELAY = 4'b0000;
defparam \cam_pclk~input .OUT_DELAY = 1'b0;
defparam \cam_pclk~input .IN_DATA_DELAY = 3'b000;
defparam \cam_pclk~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_pdown~output (
	.padio(cam_pdown),
	.datain(gnd),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \cam_pdown~output .coord_x = 22;
defparam \cam_pdown~output .coord_y = 0;
defparam \cam_pdown~output .coord_z = 0;
defparam \cam_pdown~output .IN_ASYNC_MODE = 1'b0;
defparam \cam_pdown~output .IN_SYNC_MODE = 1'b0;
defparam \cam_pdown~output .IN_POWERUP = 1'b0;
defparam \cam_pdown~output .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_pdown~output .IN_SYNC_DISABLE = 1'b0;
defparam \cam_pdown~output .OUT_REG_MODE = 1'b0;
defparam \cam_pdown~output .OUT_ASYNC_MODE = 1'b0;
defparam \cam_pdown~output .OUT_SYNC_MODE = 1'b0;
defparam \cam_pdown~output .OUT_POWERUP = 1'b0;
defparam \cam_pdown~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_pdown~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_pdown~output .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_pdown~output .OUT_DDIO = 1'b0;
defparam \cam_pdown~output .OE_REG_MODE = 1'b0;
defparam \cam_pdown~output .OE_ASYNC_MODE = 1'b0;
defparam \cam_pdown~output .OE_SYNC_MODE = 1'b0;
defparam \cam_pdown~output .OE_POWERUP = 1'b0;
defparam \cam_pdown~output .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_pdown~output .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_pdown~output .OE_SYNC_DISABLE = 1'b0;
defparam \cam_pdown~output .OE_DDIO = 1'b0;
defparam \cam_pdown~output .CFG_TRI_INPUT = 1'b0;
defparam \cam_pdown~output .CFG_PULL_UP = 1'b0;
defparam \cam_pdown~output .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_pdown~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_pdown~output .CFG_PDRV = 7'b0011010;
defparam \cam_pdown~output .CFG_NDRV = 7'b0011000;
defparam \cam_pdown~output .CFG_KEEP = 2'b00;
defparam \cam_pdown~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_pdown~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_pdown~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_pdown~output .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_pdown~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_pdown~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_pdown~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_pdown~output .CFG_OSCDIV = 2'b00;
defparam \cam_pdown~output .CFG_ROCTUSR = 1'b0;
defparam \cam_pdown~output .CFG_SEL_CUA = 1'b0;
defparam \cam_pdown~output .CFG_ROCT_EN = 1'b0;
defparam \cam_pdown~output .INPUT_ONLY = 1'b0;
defparam \cam_pdown~output .DPCLK_DELAY = 4'b0000;
defparam \cam_pdown~output .OUT_DELAY = 1'b0;
defparam \cam_pdown~output .IN_DATA_DELAY = 3'b000;
defparam \cam_pdown~output .IN_REG_DELAY = 3'b000;

alta_dio \cam_reset~output (
	.padio(cam_reset),
	.datain(!\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \cam_reset~output .coord_x = 22;
defparam \cam_reset~output .coord_y = 0;
defparam \cam_reset~output .coord_z = 1;
defparam \cam_reset~output .IN_ASYNC_MODE = 1'b0;
defparam \cam_reset~output .IN_SYNC_MODE = 1'b0;
defparam \cam_reset~output .IN_POWERUP = 1'b0;
defparam \cam_reset~output .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_reset~output .IN_SYNC_DISABLE = 1'b0;
defparam \cam_reset~output .OUT_REG_MODE = 1'b0;
defparam \cam_reset~output .OUT_ASYNC_MODE = 1'b0;
defparam \cam_reset~output .OUT_SYNC_MODE = 1'b0;
defparam \cam_reset~output .OUT_POWERUP = 1'b0;
defparam \cam_reset~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_reset~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_reset~output .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_reset~output .OUT_DDIO = 1'b0;
defparam \cam_reset~output .OE_REG_MODE = 1'b0;
defparam \cam_reset~output .OE_ASYNC_MODE = 1'b0;
defparam \cam_reset~output .OE_SYNC_MODE = 1'b0;
defparam \cam_reset~output .OE_POWERUP = 1'b0;
defparam \cam_reset~output .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_reset~output .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_reset~output .OE_SYNC_DISABLE = 1'b0;
defparam \cam_reset~output .OE_DDIO = 1'b0;
defparam \cam_reset~output .CFG_TRI_INPUT = 1'b0;
defparam \cam_reset~output .CFG_PULL_UP = 1'b0;
defparam \cam_reset~output .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_reset~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_reset~output .CFG_PDRV = 7'b0011010;
defparam \cam_reset~output .CFG_NDRV = 7'b0011000;
defparam \cam_reset~output .CFG_KEEP = 2'b00;
defparam \cam_reset~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_reset~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_reset~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_reset~output .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_reset~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_reset~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_reset~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_reset~output .CFG_OSCDIV = 2'b00;
defparam \cam_reset~output .CFG_ROCTUSR = 1'b0;
defparam \cam_reset~output .CFG_SEL_CUA = 1'b0;
defparam \cam_reset~output .CFG_ROCT_EN = 1'b0;
defparam \cam_reset~output .INPUT_ONLY = 1'b0;
defparam \cam_reset~output .DPCLK_DELAY = 4'b0000;
defparam \cam_reset~output .OUT_DELAY = 1'b0;
defparam \cam_reset~output .IN_DATA_DELAY = 3'b000;
defparam \cam_reset~output .IN_REG_DELAY = 3'b000;

alta_dio \cam_scl~output (
	.padio(cam_scl),
	.datain(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10_combout ),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \cam_scl~output .coord_x = 0;
defparam \cam_scl~output .coord_y = 13;
defparam \cam_scl~output .coord_z = 2;
defparam \cam_scl~output .IN_ASYNC_MODE = 1'b0;
defparam \cam_scl~output .IN_SYNC_MODE = 1'b0;
defparam \cam_scl~output .IN_POWERUP = 1'b0;
defparam \cam_scl~output .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_scl~output .IN_SYNC_DISABLE = 1'b0;
defparam \cam_scl~output .OUT_REG_MODE = 1'b0;
defparam \cam_scl~output .OUT_ASYNC_MODE = 1'b0;
defparam \cam_scl~output .OUT_SYNC_MODE = 1'b0;
defparam \cam_scl~output .OUT_POWERUP = 1'b0;
defparam \cam_scl~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_scl~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_scl~output .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_scl~output .OUT_DDIO = 1'b0;
defparam \cam_scl~output .OE_REG_MODE = 1'b0;
defparam \cam_scl~output .OE_ASYNC_MODE = 1'b0;
defparam \cam_scl~output .OE_SYNC_MODE = 1'b0;
defparam \cam_scl~output .OE_POWERUP = 1'b0;
defparam \cam_scl~output .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_scl~output .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_scl~output .OE_SYNC_DISABLE = 1'b0;
defparam \cam_scl~output .OE_DDIO = 1'b0;
defparam \cam_scl~output .CFG_TRI_INPUT = 1'b0;
defparam \cam_scl~output .CFG_PULL_UP = 1'b0;
defparam \cam_scl~output .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_scl~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_scl~output .CFG_PDRV = 7'b0011010;
defparam \cam_scl~output .CFG_NDRV = 7'b0011000;
defparam \cam_scl~output .CFG_KEEP = 2'b00;
defparam \cam_scl~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_scl~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_scl~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_scl~output .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_scl~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_scl~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_scl~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_scl~output .CFG_OSCDIV = 2'b00;
defparam \cam_scl~output .CFG_ROCTUSR = 1'b0;
defparam \cam_scl~output .CFG_SEL_CUA = 1'b0;
defparam \cam_scl~output .CFG_ROCT_EN = 1'b0;
defparam \cam_scl~output .INPUT_ONLY = 1'b0;
defparam \cam_scl~output .DPCLK_DELAY = 4'b0000;
defparam \cam_scl~output .OUT_DELAY = 1'b0;
defparam \cam_scl~output .IN_DATA_DELAY = 3'b000;
defparam \cam_scl~output .IN_REG_DELAY = 3'b000;

alta_dio \cam_sda~output (
	.padio(cam_sda),
	.datain(!\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.datainh(gnd),
	.oe(\camera_if_inst|u_I2C_AV_Config|u0|SDO~4_combout ),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_sda~input_o ),
	.regout());
defparam \cam_sda~output .coord_x = 0;
defparam \cam_sda~output .coord_y = 13;
defparam \cam_sda~output .coord_z = 1;
defparam \cam_sda~output .IN_ASYNC_MODE = 1'b0;
defparam \cam_sda~output .IN_SYNC_MODE = 1'b0;
defparam \cam_sda~output .IN_POWERUP = 1'b0;
defparam \cam_sda~output .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_sda~output .IN_SYNC_DISABLE = 1'b0;
defparam \cam_sda~output .OUT_REG_MODE = 1'b0;
defparam \cam_sda~output .OUT_ASYNC_MODE = 1'b0;
defparam \cam_sda~output .OUT_SYNC_MODE = 1'b0;
defparam \cam_sda~output .OUT_POWERUP = 1'b0;
defparam \cam_sda~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_sda~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_sda~output .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_sda~output .OUT_DDIO = 1'b0;
defparam \cam_sda~output .OE_REG_MODE = 1'b0;
defparam \cam_sda~output .OE_ASYNC_MODE = 1'b0;
defparam \cam_sda~output .OE_SYNC_MODE = 1'b0;
defparam \cam_sda~output .OE_POWERUP = 1'b0;
defparam \cam_sda~output .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_sda~output .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_sda~output .OE_SYNC_DISABLE = 1'b0;
defparam \cam_sda~output .OE_DDIO = 1'b0;
defparam \cam_sda~output .CFG_TRI_INPUT = 1'b0;
defparam \cam_sda~output .CFG_PULL_UP = 1'b0;
defparam \cam_sda~output .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_sda~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_sda~output .CFG_PDRV = 7'b0011010;
defparam \cam_sda~output .CFG_NDRV = 7'b0011000;
defparam \cam_sda~output .CFG_KEEP = 2'b00;
defparam \cam_sda~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_sda~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_sda~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_sda~output .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_sda~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_sda~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_sda~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_sda~output .CFG_OSCDIV = 2'b00;
defparam \cam_sda~output .CFG_ROCTUSR = 1'b0;
defparam \cam_sda~output .CFG_SEL_CUA = 1'b0;
defparam \cam_sda~output .CFG_ROCT_EN = 1'b0;
defparam \cam_sda~output .INPUT_ONLY = 1'b0;
defparam \cam_sda~output .DPCLK_DELAY = 4'b0000;
defparam \cam_sda~output .OUT_DELAY = 1'b0;
defparam \cam_sda~output .IN_DATA_DELAY = 3'b000;
defparam \cam_sda~output .IN_REG_DELAY = 3'b000;

alta_dio \cam_vsync~input (
	.padio(cam_vsync),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_vsync~input_o ),
	.regout());
defparam \cam_vsync~input .coord_x = 0;
defparam \cam_vsync~input .coord_y = 9;
defparam \cam_vsync~input .coord_z = 2;
defparam \cam_vsync~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_vsync~input .IN_SYNC_MODE = 1'b0;
defparam \cam_vsync~input .IN_POWERUP = 1'b0;
defparam \cam_vsync~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_vsync~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_vsync~input .OUT_REG_MODE = 1'b0;
defparam \cam_vsync~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_vsync~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_vsync~input .OUT_POWERUP = 1'b0;
defparam \cam_vsync~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_vsync~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_vsync~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_vsync~input .OUT_DDIO = 1'b0;
defparam \cam_vsync~input .OE_REG_MODE = 1'b0;
defparam \cam_vsync~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_vsync~input .OE_SYNC_MODE = 1'b0;
defparam \cam_vsync~input .OE_POWERUP = 1'b0;
defparam \cam_vsync~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_vsync~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_vsync~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_vsync~input .OE_DDIO = 1'b0;
defparam \cam_vsync~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_vsync~input .CFG_PULL_UP = 1'b0;
defparam \cam_vsync~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_vsync~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_vsync~input .CFG_PDRV = 7'b0011010;
defparam \cam_vsync~input .CFG_NDRV = 7'b0011000;
defparam \cam_vsync~input .CFG_KEEP = 2'b00;
defparam \cam_vsync~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_vsync~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_vsync~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_vsync~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_vsync~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_vsync~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_vsync~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_vsync~input .CFG_OSCDIV = 2'b00;
defparam \cam_vsync~input .CFG_ROCTUSR = 1'b0;
defparam \cam_vsync~input .CFG_SEL_CUA = 1'b0;
defparam \cam_vsync~input .CFG_ROCT_EN = 1'b0;
defparam \cam_vsync~input .INPUT_ONLY = 1'b0;
defparam \cam_vsync~input .DPCLK_DELAY = 4'b0000;
defparam \cam_vsync~input .OUT_DELAY = 1'b0;
defparam \cam_vsync~input .IN_DATA_DELAY = 3'b000;
defparam \cam_vsync~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_xclk~output (
	.padio(cam_xclk),
	.datain(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \cam_xclk~output .coord_x = 0;
defparam \cam_xclk~output .coord_y = 5;
defparam \cam_xclk~output .coord_z = 0;
defparam \cam_xclk~output .IN_ASYNC_MODE = 1'b0;
defparam \cam_xclk~output .IN_SYNC_MODE = 1'b0;
defparam \cam_xclk~output .IN_POWERUP = 1'b0;
defparam \cam_xclk~output .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_xclk~output .IN_SYNC_DISABLE = 1'b0;
defparam \cam_xclk~output .OUT_REG_MODE = 1'b0;
defparam \cam_xclk~output .OUT_ASYNC_MODE = 1'b0;
defparam \cam_xclk~output .OUT_SYNC_MODE = 1'b0;
defparam \cam_xclk~output .OUT_POWERUP = 1'b0;
defparam \cam_xclk~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_xclk~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_xclk~output .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_xclk~output .OUT_DDIO = 1'b0;
defparam \cam_xclk~output .OE_REG_MODE = 1'b0;
defparam \cam_xclk~output .OE_ASYNC_MODE = 1'b0;
defparam \cam_xclk~output .OE_SYNC_MODE = 1'b0;
defparam \cam_xclk~output .OE_POWERUP = 1'b0;
defparam \cam_xclk~output .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_xclk~output .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_xclk~output .OE_SYNC_DISABLE = 1'b0;
defparam \cam_xclk~output .OE_DDIO = 1'b0;
defparam \cam_xclk~output .CFG_TRI_INPUT = 1'b0;
defparam \cam_xclk~output .CFG_PULL_UP = 1'b0;
defparam \cam_xclk~output .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_xclk~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_xclk~output .CFG_PDRV = 7'b0011010;
defparam \cam_xclk~output .CFG_NDRV = 7'b0011000;
defparam \cam_xclk~output .CFG_KEEP = 2'b00;
defparam \cam_xclk~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_xclk~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_xclk~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_xclk~output .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_xclk~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_xclk~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_xclk~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_xclk~output .CFG_OSCDIV = 2'b00;
defparam \cam_xclk~output .CFG_ROCTUSR = 1'b0;
defparam \cam_xclk~output .CFG_SEL_CUA = 1'b0;
defparam \cam_xclk~output .CFG_ROCT_EN = 1'b0;
defparam \cam_xclk~output .INPUT_ONLY = 1'b0;
defparam \cam_xclk~output .DPCLK_DELAY = 4'b0000;
defparam \cam_xclk~output .OUT_DELAY = 1'b0;
defparam \cam_xclk~output .IN_DATA_DELAY = 3'b000;
defparam \cam_xclk~output .IN_REG_DELAY = 3'b000;

alta_slice \camera_if_inst|Equal0~0 (
	.A(\camera_if_inst|v_cnt [1]),
	.B(\camera_if_inst|v_cnt [3]),
	.C(\camera_if_inst|v_cnt [2]),
	.D(\camera_if_inst|v_cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal0~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal0~0 .coord_x = 12;
defparam \camera_if_inst|Equal0~0 .coord_y = 16;
defparam \camera_if_inst|Equal0~0 .coord_z = 1;
defparam \camera_if_inst|Equal0~0 .mask = 16'hFFFE;
defparam \camera_if_inst|Equal0~0 .modeMux = 1'b0;
defparam \camera_if_inst|Equal0~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal0~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal0~0 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal0~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal0~1 (
	.A(\camera_if_inst|v_cnt [5]),
	.B(\camera_if_inst|v_cnt [6]),
	.C(\camera_if_inst|v_cnt [7]),
	.D(\camera_if_inst|v_cnt [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal0~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal0~1 .coord_x = 12;
defparam \camera_if_inst|Equal0~1 .coord_y = 16;
defparam \camera_if_inst|Equal0~1 .coord_z = 4;
defparam \camera_if_inst|Equal0~1 .mask = 16'hFFFE;
defparam \camera_if_inst|Equal0~1 .modeMux = 1'b0;
defparam \camera_if_inst|Equal0~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal0~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal0~1 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal0~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal0~2 (
	.A(\camera_if_inst|v_cnt [8]),
	.B(\camera_if_inst|v_cnt [10]),
	.C(\camera_if_inst|v_cnt [9]),
	.D(\camera_if_inst|v_cnt [11]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal0~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal0~2 .coord_x = 12;
defparam \camera_if_inst|Equal0~2 .coord_y = 16;
defparam \camera_if_inst|Equal0~2 .coord_z = 6;
defparam \camera_if_inst|Equal0~2 .mask = 16'hFFFE;
defparam \camera_if_inst|Equal0~2 .modeMux = 1'b0;
defparam \camera_if_inst|Equal0~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal0~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal0~2 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal0~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal0~3 (
	.A(\camera_if_inst|v_cnt [14]),
	.B(\camera_if_inst|v_cnt [12]),
	.C(\camera_if_inst|v_cnt [13]),
	.D(\camera_if_inst|v_cnt [15]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal0~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal0~3 .coord_x = 12;
defparam \camera_if_inst|Equal0~3 .coord_y = 16;
defparam \camera_if_inst|Equal0~3 .coord_z = 3;
defparam \camera_if_inst|Equal0~3 .mask = 16'hFFFE;
defparam \camera_if_inst|Equal0~3 .modeMux = 1'b0;
defparam \camera_if_inst|Equal0~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal0~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal0~3 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal0~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal0~4 (
	.A(\camera_if_inst|Equal0~3_combout ),
	.B(\camera_if_inst|Equal0~1_combout ),
	.C(\camera_if_inst|Equal0~0_combout ),
	.D(\camera_if_inst|Equal0~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal0~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal0~4 .coord_x = 12;
defparam \camera_if_inst|Equal0~4 .coord_y = 16;
defparam \camera_if_inst|Equal0~4 .coord_z = 0;
defparam \camera_if_inst|Equal0~4 .mask = 16'hFFFE;
defparam \camera_if_inst|Equal0~4 .modeMux = 1'b0;
defparam \camera_if_inst|Equal0~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal0~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal0~4 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal0~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal2~0 (
	.A(\camera_if_inst|f_cnt [2]),
	.B(\camera_if_inst|f_cnt [1]),
	.C(vcc),
	.D(\camera_if_inst|f_cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal2~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal2~0 .coord_x = 8;
defparam \camera_if_inst|Equal2~0 .coord_y = 12;
defparam \camera_if_inst|Equal2~0 .coord_z = 9;
defparam \camera_if_inst|Equal2~0 .mask = 16'h8800;
defparam \camera_if_inst|Equal2~0 .modeMux = 1'b0;
defparam \camera_if_inst|Equal2~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal2~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal2~0 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal2~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal3~0 (
	.A(vcc),
	.B(vcc),
	.C(\camera_if_inst|h_cnt [0]),
	.D(\camera_if_inst|h_cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal3~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal3~0 .coord_x = 8;
defparam \camera_if_inst|Equal3~0 .coord_y = 12;
defparam \camera_if_inst|Equal3~0 .coord_z = 0;
defparam \camera_if_inst|Equal3~0 .mask = 16'h0FFF;
defparam \camera_if_inst|Equal3~0 .modeMux = 1'b0;
defparam \camera_if_inst|Equal3~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal3~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal3~0 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal3~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal3~1 (
	.A(\camera_if_inst|h_cnt [4]),
	.B(\camera_if_inst|h_cnt [6]),
	.C(\camera_if_inst|h_cnt [7]),
	.D(\camera_if_inst|h_cnt [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal3~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal3~1 .coord_x = 8;
defparam \camera_if_inst|Equal3~1 .coord_y = 12;
defparam \camera_if_inst|Equal3~1 .coord_z = 2;
defparam \camera_if_inst|Equal3~1 .mask = 16'hF7FF;
defparam \camera_if_inst|Equal3~1 .modeMux = 1'b0;
defparam \camera_if_inst|Equal3~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal3~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal3~1 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal3~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal3~2 (
	.A(\camera_if_inst|Equal3~0_combout ),
	.B(\camera_if_inst|Equal3~1_combout ),
	.C(\camera_if_inst|h_cnt [2]),
	.D(\camera_if_inst|h_cnt [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal3~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal3~2 .coord_x = 8;
defparam \camera_if_inst|Equal3~2 .coord_y = 12;
defparam \camera_if_inst|Equal3~2 .coord_z = 15;
defparam \camera_if_inst|Equal3~2 .mask = 16'hEFFF;
defparam \camera_if_inst|Equal3~2 .modeMux = 1'b0;
defparam \camera_if_inst|Equal3~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal3~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal3~2 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal3~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal3~3 (
	.A(\camera_if_inst|h_cnt [9]),
	.B(\camera_if_inst|h_cnt [11]),
	.C(\camera_if_inst|h_cnt [10]),
	.D(\camera_if_inst|h_cnt [8]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal3~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal3~3 .coord_x = 8;
defparam \camera_if_inst|Equal3~3 .coord_y = 12;
defparam \camera_if_inst|Equal3~3 .coord_z = 8;
defparam \camera_if_inst|Equal3~3 .mask = 16'hFFFD;
defparam \camera_if_inst|Equal3~3 .modeMux = 1'b0;
defparam \camera_if_inst|Equal3~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal3~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal3~3 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal3~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal3~4 (
	.A(\camera_if_inst|h_cnt [15]),
	.B(\camera_if_inst|h_cnt [14]),
	.C(\camera_if_inst|h_cnt [13]),
	.D(\camera_if_inst|h_cnt [12]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal3~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal3~4 .coord_x = 8;
defparam \camera_if_inst|Equal3~4 .coord_y = 12;
defparam \camera_if_inst|Equal3~4 .coord_z = 13;
defparam \camera_if_inst|Equal3~4 .mask = 16'hFFFE;
defparam \camera_if_inst|Equal3~4 .modeMux = 1'b0;
defparam \camera_if_inst|Equal3~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal3~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal3~4 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal3~4 .CarryEnb = 1'b1;

alta_io_gclk \camera_if_inst|Equal4~0clkctrl (
	.inclk(\camera_if_inst|Equal4~0_combout ),
	.outclk(\camera_if_inst|Equal4~0clkctrl_outclk ));
defparam \camera_if_inst|Equal4~0clkctrl .coord_x = 0;
defparam \camera_if_inst|Equal4~0clkctrl .coord_y = 12;
defparam \camera_if_inst|Equal4~0clkctrl .coord_z = 4;

alta_slice \camera_if_inst|cam_data_r0[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cam_data[0]~input_o ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [0]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r0[0]~feeder_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [0]));
defparam \camera_if_inst|cam_data_r0[0] .coord_x = 17;
defparam \camera_if_inst|cam_data_r0[0] .coord_y = 12;
defparam \camera_if_inst|cam_data_r0[0] .coord_z = 11;
defparam \camera_if_inst|cam_data_r0[0] .mask = 16'hFF00;
defparam \camera_if_inst|cam_data_r0[0] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[0] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r0[0] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[1] (
	.A(),
	.B(),
	.C(\cam_data[1]~input_o ),
	.D(),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [1]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(SyncReset_X4_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X4_Y7_VCC),
	.LutOut(),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [1]));
defparam \camera_if_inst|cam_data_r0[1] .coord_x = 17;
defparam \camera_if_inst|cam_data_r0[1] .coord_y = 12;
defparam \camera_if_inst|cam_data_r0[1] .coord_z = 8;
defparam \camera_if_inst|cam_data_r0[1] .mask = 16'hFFFF;
defparam \camera_if_inst|cam_data_r0[1] .modeMux = 1'b1;
defparam \camera_if_inst|cam_data_r0[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[1] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_data_r0[1] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[2] (
	.A(),
	.B(),
	.C(\cam_data[2]~input_o ),
	.D(),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [2]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(SyncReset_X4_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X4_Y7_VCC),
	.LutOut(),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [2]));
defparam \camera_if_inst|cam_data_r0[2] .coord_x = 17;
defparam \camera_if_inst|cam_data_r0[2] .coord_y = 12;
defparam \camera_if_inst|cam_data_r0[2] .coord_z = 15;
defparam \camera_if_inst|cam_data_r0[2] .mask = 16'hFFFF;
defparam \camera_if_inst|cam_data_r0[2] .modeMux = 1'b1;
defparam \camera_if_inst|cam_data_r0[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[2] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_data_r0[2] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[3] (
	.A(\camera_if_inst|cam_data_r0 [0]),
	.B(\camera_if_inst|cam_data_r0 [1]),
	.C(\cam_data[3]~input_o ),
	.D(\camera_if_inst|cam_data_r0 [2]),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [3]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(SyncReset_X4_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X4_Y7_VCC),
	.LutOut(\camera_if_inst|Equal1~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [3]));
defparam \camera_if_inst|cam_data_r0[3] .coord_x = 17;
defparam \camera_if_inst|cam_data_r0[3] .coord_y = 12;
defparam \camera_if_inst|cam_data_r0[3] .coord_z = 3;
defparam \camera_if_inst|cam_data_r0[3] .mask = 16'hFFFE;
defparam \camera_if_inst|cam_data_r0[3] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[3] .FeedbackMux = 1'b1;
defparam \camera_if_inst|cam_data_r0[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[3] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_data_r0[3] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[4] (
	.A(),
	.B(),
	.C(\cam_data[4]~input_o ),
	.D(),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [4]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(SyncReset_X4_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X4_Y7_VCC),
	.LutOut(),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [4]));
defparam \camera_if_inst|cam_data_r0[4] .coord_x = 17;
defparam \camera_if_inst|cam_data_r0[4] .coord_y = 12;
defparam \camera_if_inst|cam_data_r0[4] .coord_z = 9;
defparam \camera_if_inst|cam_data_r0[4] .mask = 16'hFFFF;
defparam \camera_if_inst|cam_data_r0[4] .modeMux = 1'b1;
defparam \camera_if_inst|cam_data_r0[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[4] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_data_r0[4] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cam_data[5]~input_o ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [5]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r0[5]~feeder_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [5]));
defparam \camera_if_inst|cam_data_r0[5] .coord_x = 17;
defparam \camera_if_inst|cam_data_r0[5] .coord_y = 12;
defparam \camera_if_inst|cam_data_r0[5] .coord_z = 1;
defparam \camera_if_inst|cam_data_r0[5] .mask = 16'hFF00;
defparam \camera_if_inst|cam_data_r0[5] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[5] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[5] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r0[5] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[6] (
	.A(),
	.B(),
	.C(\cam_data[6]~input_o ),
	.D(),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [6]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(SyncReset_X4_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X4_Y7_VCC),
	.LutOut(),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [6]));
defparam \camera_if_inst|cam_data_r0[6] .coord_x = 17;
defparam \camera_if_inst|cam_data_r0[6] .coord_y = 12;
defparam \camera_if_inst|cam_data_r0[6] .coord_z = 14;
defparam \camera_if_inst|cam_data_r0[6] .mask = 16'hFFFF;
defparam \camera_if_inst|cam_data_r0[6] .modeMux = 1'b1;
defparam \camera_if_inst|cam_data_r0[6] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[6] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[6] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_data_r0[6] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[7] (
	.A(\camera_if_inst|cam_data_r0 [5]),
	.B(\camera_if_inst|cam_data_r0 [6]),
	.C(\cam_data[7]~input_o ),
	.D(\camera_if_inst|cam_data_r0 [4]),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [7]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(SyncReset_X4_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X4_Y7_VCC),
	.LutOut(\camera_if_inst|Equal1~1_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [7]));
defparam \camera_if_inst|cam_data_r0[7] .coord_x = 17;
defparam \camera_if_inst|cam_data_r0[7] .coord_y = 12;
defparam \camera_if_inst|cam_data_r0[7] .coord_z = 7;
defparam \camera_if_inst|cam_data_r0[7] .mask = 16'hFFFE;
defparam \camera_if_inst|cam_data_r0[7] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[7] .FeedbackMux = 1'b1;
defparam \camera_if_inst|cam_data_r0[7] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[7] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_data_r0[7] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[0] (
	.A(\camera_if_inst|cam_data_r0 [0]),
	.B(\camera_if_inst|Equal0~4_combout ),
	.C(\camera_if_inst|Equal1~1_combout ),
	.D(\camera_if_inst|Equal1~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [0]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [0]));
defparam \camera_if_inst|cam_data_r1[0] .coord_x = 17;
defparam \camera_if_inst|cam_data_r1[0] .coord_y = 12;
defparam \camera_if_inst|cam_data_r1[0] .coord_z = 10;
defparam \camera_if_inst|cam_data_r1[0] .mask = 16'h888C;
defparam \camera_if_inst|cam_data_r1[0] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[0] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[0] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[1] (
	.A(\camera_if_inst|Equal0~4_combout ),
	.B(\camera_if_inst|cam_data_r0 [1]),
	.C(\camera_if_inst|Equal1~1_combout ),
	.D(\camera_if_inst|Equal1~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [1]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~7_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [1]));
defparam \camera_if_inst|cam_data_r1[1] .coord_x = 17;
defparam \camera_if_inst|cam_data_r1[1] .coord_y = 12;
defparam \camera_if_inst|cam_data_r1[1] .coord_z = 5;
defparam \camera_if_inst|cam_data_r1[1] .mask = 16'h8880;
defparam \camera_if_inst|cam_data_r1[1] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[1] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[1] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[2] (
	.A(\camera_if_inst|Equal0~4_combout ),
	.B(\camera_if_inst|cam_data_r0 [2]),
	.C(\camera_if_inst|Equal1~1_combout ),
	.D(\camera_if_inst|Equal1~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [2]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~1_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [2]));
defparam \camera_if_inst|cam_data_r1[2] .coord_x = 17;
defparam \camera_if_inst|cam_data_r1[2] .coord_y = 12;
defparam \camera_if_inst|cam_data_r1[2] .coord_z = 12;
defparam \camera_if_inst|cam_data_r1[2] .mask = 16'h8880;
defparam \camera_if_inst|cam_data_r1[2] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[2] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[2] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[3] (
	.A(\camera_if_inst|cam_data_r0 [3]),
	.B(\camera_if_inst|Equal0~4_combout ),
	.C(\camera_if_inst|Equal1~1_combout ),
	.D(\camera_if_inst|Equal1~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [3]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~5_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [3]));
defparam \camera_if_inst|cam_data_r1[3] .coord_x = 17;
defparam \camera_if_inst|cam_data_r1[3] .coord_y = 12;
defparam \camera_if_inst|cam_data_r1[3] .coord_z = 6;
defparam \camera_if_inst|cam_data_r1[3] .mask = 16'h8880;
defparam \camera_if_inst|cam_data_r1[3] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[3] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[3] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[3] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[4] (
	.A(\camera_if_inst|cam_data_r0 [4]),
	.B(\camera_if_inst|Equal0~4_combout ),
	.C(\camera_if_inst|Equal1~1_combout ),
	.D(\camera_if_inst|Equal1~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [4]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~3_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [4]));
defparam \camera_if_inst|cam_data_r1[4] .coord_x = 17;
defparam \camera_if_inst|cam_data_r1[4] .coord_y = 12;
defparam \camera_if_inst|cam_data_r1[4] .coord_z = 13;
defparam \camera_if_inst|cam_data_r1[4] .mask = 16'h8880;
defparam \camera_if_inst|cam_data_r1[4] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[4] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[4] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[5] (
	.A(\camera_if_inst|cam_data_r0 [5]),
	.B(\camera_if_inst|Equal0~4_combout ),
	.C(\camera_if_inst|Equal1~1_combout ),
	.D(\camera_if_inst|Equal1~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [5]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~6_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [5]));
defparam \camera_if_inst|cam_data_r1[5] .coord_x = 17;
defparam \camera_if_inst|cam_data_r1[5] .coord_y = 12;
defparam \camera_if_inst|cam_data_r1[5] .coord_z = 4;
defparam \camera_if_inst|cam_data_r1[5] .mask = 16'h8880;
defparam \camera_if_inst|cam_data_r1[5] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[5] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[5] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[5] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[6] (
	.A(\camera_if_inst|Equal1~0_combout ),
	.B(\camera_if_inst|cam_data_r0 [6]),
	.C(\camera_if_inst|Equal1~1_combout ),
	.D(\camera_if_inst|Equal0~4_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [6]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [6]));
defparam \camera_if_inst|cam_data_r1[6] .coord_x = 17;
defparam \camera_if_inst|cam_data_r1[6] .coord_y = 12;
defparam \camera_if_inst|cam_data_r1[6] .coord_z = 2;
defparam \camera_if_inst|cam_data_r1[6] .mask = 16'hC800;
defparam \camera_if_inst|cam_data_r1[6] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[6] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[6] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[6] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[6] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[7] (
	.A(\camera_if_inst|cam_data_r0 [7]),
	.B(\camera_if_inst|Equal0~4_combout ),
	.C(\camera_if_inst|Equal1~1_combout ),
	.D(\camera_if_inst|Equal1~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [7]),
	.Clk(\cam_pclk~input_o_X4_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X4_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~4_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [7]));
defparam \camera_if_inst|cam_data_r1[7] .coord_x = 17;
defparam \camera_if_inst|cam_data_r1[7] .coord_y = 12;
defparam \camera_if_inst|cam_data_r1[7] .coord_z = 0;
defparam \camera_if_inst|cam_data_r1[7] .mask = 16'h8880;
defparam \camera_if_inst|cam_data_r1[7] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[7] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[7] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[7] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[7] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_hsync_r[0] (
	.A(vcc),
	.B(\camera_if_inst|f_cnt [3]),
	.C(\cam_hsync~input_o ),
	.D(\camera_if_inst|Equal2~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_hsync_r [0]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_hsync_r~1_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_hsync_r [0]));
defparam \camera_if_inst|cam_hsync_r[0] .coord_x = 8;
defparam \camera_if_inst|cam_hsync_r[0] .coord_y = 12;
defparam \camera_if_inst|cam_hsync_r[0] .coord_z = 3;
defparam \camera_if_inst|cam_hsync_r[0] .mask = 16'hC000;
defparam \camera_if_inst|cam_hsync_r[0] .modeMux = 1'b0;
defparam \camera_if_inst|cam_hsync_r[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_hsync_r[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_hsync_r[0] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_hsync_r[0] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_hsync_r[1] (
	.A(\camera_if_inst|cam_hsync_r [0]),
	.B(\camera_if_inst|f_cnt [3]),
	.C(vcc),
	.D(\camera_if_inst|Equal2~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_hsync_r [1]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_hsync_r~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_hsync_r [1]));
defparam \camera_if_inst|cam_hsync_r[1] .coord_x = 8;
defparam \camera_if_inst|cam_hsync_r[1] .coord_y = 12;
defparam \camera_if_inst|cam_hsync_r[1] .coord_z = 4;
defparam \camera_if_inst|cam_hsync_r[1] .mask = 16'h8800;
defparam \camera_if_inst|cam_hsync_r[1] .modeMux = 1'b0;
defparam \camera_if_inst|cam_hsync_r[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_hsync_r[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_hsync_r[1] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_hsync_r[1] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_vsync_r[0] (
	.A(\camera_if_inst|cam_vsync_r [1]),
	.B(\camera_if_inst|f_cnt [3]),
	.C(\cam_vsync~input_o ),
	.D(\camera_if_inst|Equal2~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_vsync_r [0]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(SyncReset_X1_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_VCC),
	.LutOut(\camera_if_inst|f_cnt[3]~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_vsync_r [0]));
defparam \camera_if_inst|cam_vsync_r[0] .coord_x = 8;
defparam \camera_if_inst|cam_vsync_r[0] .coord_y = 12;
defparam \camera_if_inst|cam_vsync_r[0] .coord_z = 10;
defparam \camera_if_inst|cam_vsync_r[0] .mask = 16'h020A;
defparam \camera_if_inst|cam_vsync_r[0] .modeMux = 1'b0;
defparam \camera_if_inst|cam_vsync_r[0] .FeedbackMux = 1'b1;
defparam \camera_if_inst|cam_vsync_r[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_vsync_r[0] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_vsync_r[0] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_vsync_r[1] (
	.A(vcc),
	.B(\camera_if_inst|cam_vsync_r [0]),
	.C(\camera_if_inst|cam_vsync_r [0]),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|cam_vsync_r [1]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(SyncReset_X1_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_VCC),
	.LutOut(\camera_if_inst|Equal4~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_vsync_r [1]));
defparam \camera_if_inst|cam_vsync_r[1] .coord_x = 8;
defparam \camera_if_inst|cam_vsync_r[1] .coord_y = 12;
defparam \camera_if_inst|cam_vsync_r[1] .coord_z = 5;
defparam \camera_if_inst|cam_vsync_r[1] .mask = 16'h3030;
defparam \camera_if_inst|cam_vsync_r[1] .modeMux = 1'b0;
defparam \camera_if_inst|cam_vsync_r[1] .FeedbackMux = 1'b1;
defparam \camera_if_inst|cam_vsync_r[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_vsync_r[1] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_vsync_r[1] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|f_cnt[0] (
	.A(\camera_if_inst|Equal4~0_combout ),
	.B(\camera_if_inst|f_cnt [3]),
	.C(vcc),
	.D(\camera_if_inst|Equal2~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|f_cnt [0]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|f_cnt[0]~5_combout ),
	.Cout(),
	.Q(\camera_if_inst|f_cnt [0]));
defparam \camera_if_inst|f_cnt[0] .coord_x = 8;
defparam \camera_if_inst|f_cnt[0] .coord_y = 12;
defparam \camera_if_inst|f_cnt[0] .coord_z = 11;
defparam \camera_if_inst|f_cnt[0] .mask = 16'hD25A;
defparam \camera_if_inst|f_cnt[0] .modeMux = 1'b0;
defparam \camera_if_inst|f_cnt[0] .FeedbackMux = 1'b1;
defparam \camera_if_inst|f_cnt[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|f_cnt[0] .BypassEn = 1'b0;
defparam \camera_if_inst|f_cnt[0] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|f_cnt[1] (
	.A(\camera_if_inst|f_cnt [0]),
	.B(vcc),
	.C(vcc),
	.D(\camera_if_inst|f_cnt[3]~2_combout ),
	.Cin(),
	.Qin(\camera_if_inst|f_cnt [1]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|f_cnt[1]~4_combout ),
	.Cout(),
	.Q(\camera_if_inst|f_cnt [1]));
defparam \camera_if_inst|f_cnt[1] .coord_x = 8;
defparam \camera_if_inst|f_cnt[1] .coord_y = 12;
defparam \camera_if_inst|f_cnt[1] .coord_z = 12;
defparam \camera_if_inst|f_cnt[1] .mask = 16'h5AF0;
defparam \camera_if_inst|f_cnt[1] .modeMux = 1'b0;
defparam \camera_if_inst|f_cnt[1] .FeedbackMux = 1'b1;
defparam \camera_if_inst|f_cnt[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|f_cnt[1] .BypassEn = 1'b0;
defparam \camera_if_inst|f_cnt[1] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|f_cnt[2] (
	.A(\camera_if_inst|f_cnt [0]),
	.B(\camera_if_inst|f_cnt [1]),
	.C(vcc),
	.D(\camera_if_inst|f_cnt[3]~2_combout ),
	.Cin(),
	.Qin(\camera_if_inst|f_cnt [2]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|f_cnt[2]~3_combout ),
	.Cout(),
	.Q(\camera_if_inst|f_cnt [2]));
defparam \camera_if_inst|f_cnt[2] .coord_x = 8;
defparam \camera_if_inst|f_cnt[2] .coord_y = 12;
defparam \camera_if_inst|f_cnt[2] .coord_z = 1;
defparam \camera_if_inst|f_cnt[2] .mask = 16'h78F0;
defparam \camera_if_inst|f_cnt[2] .modeMux = 1'b0;
defparam \camera_if_inst|f_cnt[2] .FeedbackMux = 1'b1;
defparam \camera_if_inst|f_cnt[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|f_cnt[2] .BypassEn = 1'b0;
defparam \camera_if_inst|f_cnt[2] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|f_cnt[3] (
	.A(\camera_if_inst|cam_vsync_r [1]),
	.B(\camera_if_inst|cam_vsync_r [0]),
	.C(vcc),
	.D(\camera_if_inst|Equal2~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|f_cnt [3]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|f_cnt[3]~6_combout ),
	.Cout(),
	.Q(\camera_if_inst|f_cnt [3]));
defparam \camera_if_inst|f_cnt[3] .coord_x = 8;
defparam \camera_if_inst|f_cnt[3] .coord_y = 12;
defparam \camera_if_inst|f_cnt[3] .coord_z = 7;
defparam \camera_if_inst|f_cnt[3] .mask = 16'hF2F0;
defparam \camera_if_inst|f_cnt[3] .modeMux = 1'b0;
defparam \camera_if_inst|f_cnt[3] .FeedbackMux = 1'b1;
defparam \camera_if_inst|f_cnt[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|f_cnt[3] .BypassEn = 1'b0;
defparam \camera_if_inst|f_cnt[3] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|h_cnt[0] (
	.A(\camera_if_inst|h_cnt [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|h_cnt [0]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[0]~16_combout ),
	.Cout(\camera_if_inst|h_cnt[0]~17 ),
	.Q(\camera_if_inst|h_cnt [0]));
defparam \camera_if_inst|h_cnt[0] .coord_x = 9;
defparam \camera_if_inst|h_cnt[0] .coord_y = 12;
defparam \camera_if_inst|h_cnt[0] .coord_z = 0;
defparam \camera_if_inst|h_cnt[0] .mask = 16'h55AA;
defparam \camera_if_inst|h_cnt[0] .modeMux = 1'b0;
defparam \camera_if_inst|h_cnt[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[0] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[0] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[10] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [10]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[9]~35 ),
	.Qin(\camera_if_inst|h_cnt [10]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[10]~36_combout ),
	.Cout(\camera_if_inst|h_cnt[10]~37 ),
	.Q(\camera_if_inst|h_cnt [10]));
defparam \camera_if_inst|h_cnt[10] .coord_x = 9;
defparam \camera_if_inst|h_cnt[10] .coord_y = 12;
defparam \camera_if_inst|h_cnt[10] .coord_z = 10;
defparam \camera_if_inst|h_cnt[10] .mask = 16'hC30C;
defparam \camera_if_inst|h_cnt[10] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[10] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[10] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[10] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[10] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[11] (
	.A(\camera_if_inst|h_cnt [11]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[10]~37 ),
	.Qin(\camera_if_inst|h_cnt [11]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[11]~38_combout ),
	.Cout(\camera_if_inst|h_cnt[11]~39 ),
	.Q(\camera_if_inst|h_cnt [11]));
defparam \camera_if_inst|h_cnt[11] .coord_x = 9;
defparam \camera_if_inst|h_cnt[11] .coord_y = 12;
defparam \camera_if_inst|h_cnt[11] .coord_z = 11;
defparam \camera_if_inst|h_cnt[11] .mask = 16'h5A5F;
defparam \camera_if_inst|h_cnt[11] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[11] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[11] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[11] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[11] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[12] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [12]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[11]~39 ),
	.Qin(\camera_if_inst|h_cnt [12]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[12]~40_combout ),
	.Cout(\camera_if_inst|h_cnt[12]~41 ),
	.Q(\camera_if_inst|h_cnt [12]));
defparam \camera_if_inst|h_cnt[12] .coord_x = 9;
defparam \camera_if_inst|h_cnt[12] .coord_y = 12;
defparam \camera_if_inst|h_cnt[12] .coord_z = 12;
defparam \camera_if_inst|h_cnt[12] .mask = 16'hC30C;
defparam \camera_if_inst|h_cnt[12] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[12] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[12] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[12] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[12] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[13] (
	.A(\camera_if_inst|h_cnt [13]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[12]~41 ),
	.Qin(\camera_if_inst|h_cnt [13]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[13]~42_combout ),
	.Cout(\camera_if_inst|h_cnt[13]~43 ),
	.Q(\camera_if_inst|h_cnt [13]));
defparam \camera_if_inst|h_cnt[13] .coord_x = 9;
defparam \camera_if_inst|h_cnt[13] .coord_y = 12;
defparam \camera_if_inst|h_cnt[13] .coord_z = 13;
defparam \camera_if_inst|h_cnt[13] .mask = 16'h5A5F;
defparam \camera_if_inst|h_cnt[13] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[13] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[13] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[13] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[13] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[14] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [14]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[13]~43 ),
	.Qin(\camera_if_inst|h_cnt [14]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[14]~44_combout ),
	.Cout(\camera_if_inst|h_cnt[14]~45 ),
	.Q(\camera_if_inst|h_cnt [14]));
defparam \camera_if_inst|h_cnt[14] .coord_x = 9;
defparam \camera_if_inst|h_cnt[14] .coord_y = 12;
defparam \camera_if_inst|h_cnt[14] .coord_z = 14;
defparam \camera_if_inst|h_cnt[14] .mask = 16'hC30C;
defparam \camera_if_inst|h_cnt[14] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[14] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[14] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[14] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[14] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[15] (
	.A(\camera_if_inst|h_cnt [15]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[14]~45 ),
	.Qin(\camera_if_inst|h_cnt [15]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[15]~46_combout ),
	.Cout(),
	.Q(\camera_if_inst|h_cnt [15]));
defparam \camera_if_inst|h_cnt[15] .coord_x = 9;
defparam \camera_if_inst|h_cnt[15] .coord_y = 12;
defparam \camera_if_inst|h_cnt[15] .coord_z = 15;
defparam \camera_if_inst|h_cnt[15] .mask = 16'h5A5A;
defparam \camera_if_inst|h_cnt[15] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[15] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[15] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[15] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[15] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|h_cnt[1] (
	.A(\camera_if_inst|h_cnt [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[0]~17 ),
	.Qin(\camera_if_inst|h_cnt [1]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[1]~18_combout ),
	.Cout(\camera_if_inst|h_cnt[1]~19 ),
	.Q(\camera_if_inst|h_cnt [1]));
defparam \camera_if_inst|h_cnt[1] .coord_x = 9;
defparam \camera_if_inst|h_cnt[1] .coord_y = 12;
defparam \camera_if_inst|h_cnt[1] .coord_z = 1;
defparam \camera_if_inst|h_cnt[1] .mask = 16'h5A5F;
defparam \camera_if_inst|h_cnt[1] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[1] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[1] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[2] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[1]~19 ),
	.Qin(\camera_if_inst|h_cnt [2]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[2]~20_combout ),
	.Cout(\camera_if_inst|h_cnt[2]~21 ),
	.Q(\camera_if_inst|h_cnt [2]));
defparam \camera_if_inst|h_cnt[2] .coord_x = 9;
defparam \camera_if_inst|h_cnt[2] .coord_y = 12;
defparam \camera_if_inst|h_cnt[2] .coord_z = 2;
defparam \camera_if_inst|h_cnt[2] .mask = 16'hC30C;
defparam \camera_if_inst|h_cnt[2] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[2] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[2] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[3] (
	.A(\camera_if_inst|h_cnt [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[2]~21 ),
	.Qin(\camera_if_inst|h_cnt [3]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[3]~22_combout ),
	.Cout(\camera_if_inst|h_cnt[3]~23 ),
	.Q(\camera_if_inst|h_cnt [3]));
defparam \camera_if_inst|h_cnt[3] .coord_x = 9;
defparam \camera_if_inst|h_cnt[3] .coord_y = 12;
defparam \camera_if_inst|h_cnt[3] .coord_z = 3;
defparam \camera_if_inst|h_cnt[3] .mask = 16'h5A5F;
defparam \camera_if_inst|h_cnt[3] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[3] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[3] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[3] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[4] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[3]~23 ),
	.Qin(\camera_if_inst|h_cnt [4]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[4]~24_combout ),
	.Cout(\camera_if_inst|h_cnt[4]~25 ),
	.Q(\camera_if_inst|h_cnt [4]));
defparam \camera_if_inst|h_cnt[4] .coord_x = 9;
defparam \camera_if_inst|h_cnt[4] .coord_y = 12;
defparam \camera_if_inst|h_cnt[4] .coord_z = 4;
defparam \camera_if_inst|h_cnt[4] .mask = 16'hC30C;
defparam \camera_if_inst|h_cnt[4] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[4] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[4] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[5] (
	.A(\camera_if_inst|h_cnt [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[4]~25 ),
	.Qin(\camera_if_inst|h_cnt [5]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[5]~26_combout ),
	.Cout(\camera_if_inst|h_cnt[5]~27 ),
	.Q(\camera_if_inst|h_cnt [5]));
defparam \camera_if_inst|h_cnt[5] .coord_x = 9;
defparam \camera_if_inst|h_cnt[5] .coord_y = 12;
defparam \camera_if_inst|h_cnt[5] .coord_z = 5;
defparam \camera_if_inst|h_cnt[5] .mask = 16'h5A5F;
defparam \camera_if_inst|h_cnt[5] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[5] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[5] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[5] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[6] (
	.A(\camera_if_inst|h_cnt [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[5]~27 ),
	.Qin(\camera_if_inst|h_cnt [6]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[6]~28_combout ),
	.Cout(\camera_if_inst|h_cnt[6]~29 ),
	.Q(\camera_if_inst|h_cnt [6]));
defparam \camera_if_inst|h_cnt[6] .coord_x = 9;
defparam \camera_if_inst|h_cnt[6] .coord_y = 12;
defparam \camera_if_inst|h_cnt[6] .coord_z = 6;
defparam \camera_if_inst|h_cnt[6] .mask = 16'hA50A;
defparam \camera_if_inst|h_cnt[6] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[6] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[6] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[6] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[6] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[7] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[6]~29 ),
	.Qin(\camera_if_inst|h_cnt [7]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[7]~30_combout ),
	.Cout(\camera_if_inst|h_cnt[7]~31 ),
	.Q(\camera_if_inst|h_cnt [7]));
defparam \camera_if_inst|h_cnt[7] .coord_x = 9;
defparam \camera_if_inst|h_cnt[7] .coord_y = 12;
defparam \camera_if_inst|h_cnt[7] .coord_z = 7;
defparam \camera_if_inst|h_cnt[7] .mask = 16'h3C3F;
defparam \camera_if_inst|h_cnt[7] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[7] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[7] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[7] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[7] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[8] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [8]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[7]~31 ),
	.Qin(\camera_if_inst|h_cnt [8]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[8]~32_combout ),
	.Cout(\camera_if_inst|h_cnt[8]~33 ),
	.Q(\camera_if_inst|h_cnt [8]));
defparam \camera_if_inst|h_cnt[8] .coord_x = 9;
defparam \camera_if_inst|h_cnt[8] .coord_y = 12;
defparam \camera_if_inst|h_cnt[8] .coord_z = 8;
defparam \camera_if_inst|h_cnt[8] .mask = 16'hC30C;
defparam \camera_if_inst|h_cnt[8] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[8] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[8] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[8] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[8] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[9] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [9]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[8]~33 ),
	.Qin(\camera_if_inst|h_cnt [9]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[9]~34_combout ),
	.Cout(\camera_if_inst|h_cnt[9]~35 ),
	.Q(\camera_if_inst|h_cnt [9]));
defparam \camera_if_inst|h_cnt[9] .coord_x = 9;
defparam \camera_if_inst|h_cnt[9] .coord_y = 12;
defparam \camera_if_inst|h_cnt[9] .coord_z = 9;
defparam \camera_if_inst|h_cnt[9] .mask = 16'h3C3F;
defparam \camera_if_inst|h_cnt[9] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[9] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[9] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[9] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[9] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] (
	.A(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.10~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X17_Y17_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0]~22_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .mask = 16'h78F0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .FeedbackMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1]~7_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1]~8 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .mask = 16'h6688;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1]~8 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2]~9_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2]~10 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .mask = 16'h3C3F;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2]~10 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3]~11_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3]~12 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3]~12 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4]~14_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4]~15 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4]~15 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5]~16_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5]~17 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5]~17 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6]~18_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6]~19 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6]~19 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~20_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .mask = 16'hC3C3;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 (
	.A(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.10~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|LessThan1~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .mask = 16'hA200;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan0~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [11]),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [13]),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [12]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [14]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan0~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .mask = 16'h0001;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan0~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan0~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .mask = 16'h0001;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan0~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [5]),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan0~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .mask = 16'h7F7F;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan0~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LessThan0~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [8]),
	.C(\camera_if_inst|u_I2C_AV_Config|LessThan0~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [9]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan0~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .mask = 16'h0032;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan0~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LessThan0~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LessThan0~3_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [15]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .mask = 16'h080A;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan1~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan1~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .mask = 16'h010F;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan1~1 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|LessThan1~0_combout ),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .mask = 16'hF3F3;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|Selector3~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|Selector3~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .mask = 16'h4400;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|Selector3~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|Selector3~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .mask = 16'hFFFE;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|Selector3~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|Selector3~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|Selector3~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .mask = 16'hFFFE;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X22_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~feeder_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~q ));
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .mask = 16'hAAAA;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~q ),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|i2c_en_r1~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X22_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y8_SIG ),
	.SyncReset(SyncReset_X22_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X22_Y8_VCC),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|i2c_en_r1~q ));
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .mask = 16'h3030;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .FeedbackMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [0]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0]~16_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0]~17 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [0]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .mask = 16'h55AA;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [10]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9]~35 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [10]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10]~36_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10]~37 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [10]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [11]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10]~37 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [11]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11]~38_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11]~39 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [11]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [12]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11]~39 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [12]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12]~40_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12]~41 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [12]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [13]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12]~41 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [13]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13]~42_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13]~43 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [13]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [14]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13]~43 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [14]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14]~44_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14]~45 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [14]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [15]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14]~45 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [15]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15]~46_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [15]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .mask = 16'h5A5A;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0]~17 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [1]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1]~18_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1]~19 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [1]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1]~19 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [2]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2]~20_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2]~21 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [2]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2]~21 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [3]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3]~22_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3]~23 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [3]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3]~23 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [4]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4]~24_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4]~25 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [4]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4]~25 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [5]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5]~26_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5]~27 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [5]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5]~27 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [6]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6]~28_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6]~29 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [6]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .mask = 16'hA50A;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6]~29 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [7]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7]~30_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7]~31 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [7]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .mask = 16'h3C3F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [8]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7]~31 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [8]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8]~32_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8]~33 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [8]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [9]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8]~33 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [9]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9]~34_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9]~35 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [9]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .mask = 16'h3C3F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X22_Y8_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~q ));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .mask = 16'hC3C3;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .FeedbackMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_GO (
	.A(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.00~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~1_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .mask = 16'hD500;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.B(vcc),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .mask = 16'h5500;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_WR (
	.A(\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|Selector3~2_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.00~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|Selector3~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .mask = 16'hAA08;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 (
	.A(\camera_if_inst|u_I2C_AV_Config|mSetup_ST~11_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACK~2_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.00~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mSetup_ST~12_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.00~q ));
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .mask = 16'h1050;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 (
	.A(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.10~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|LessThan1~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mSetup_ST~10_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ));
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .mask = 16'h0051;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 (
	.A(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACK~2_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.10~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mSetup_ST~13_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.10~q ));
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .mask = 16'h2000;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 (
	.A(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.00~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mSetup_ST~11_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .mask = 16'h3322;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .mask = 16'h4C00;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 (
	.A(\cam_sda~input_o ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .mask = 16'h50C0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Selector9~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .mask = 16'hCCD8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .mask = 16'h002A;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.D(\cam_sda~input_o ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .mask = 16'h1505;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|END~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Selector8~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .mask = 16'h55CD;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~3_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .mask = 16'h004C;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 (
	.A(\cam_sda~input_o ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .mask = 16'hBB33;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .mask = 16'h9000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .mask = 16'hA3B3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .mask = 16'h4500;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\cam_sda~input_o ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .mask = 16'h8A0A;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Selector9~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|END~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .mask = 16'h7745;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .mask = 16'hB000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 (
	.A(\cam_sda~input_o ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .mask = 16'hC050;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Selector8~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .mask = 16'hCCE4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .mask = 16'h4500;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\cam_sda~input_o ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .mask = 16'hA222;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|END~4_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Selector2~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .mask = 16'h5F51;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACK~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .mask = 16'h070F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACK~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .mask = 16'h4CCC;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 (
	.A(vcc),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACK~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|ACK~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACK~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .mask = 16'hFFF0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .mask = 16'h1111;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 (
	.A(vcc),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .mask = 16'h000F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .mask = 16'h1000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|END~5_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|END~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~6_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|END~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .mask = 16'hEC00;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END~0 (
	.A(vcc),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .mask = 16'hF000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .mask = 16'hA2AA;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END~2 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .mask = 16'h0033;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|END~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .mask = 16'h8000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END~4 (
	.A(vcc),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .mask = 16'hF000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|END~4_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|END~3_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|END~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .mask = 16'hECCC;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(vcc),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .mask = 16'h0055;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .mask = 16'h8000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Equal3~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .mask = 16'h0100;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Equal3~0_combout ),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Equal3~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .mask = 16'h8080;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Equal5~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .mask = 16'h2000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~29_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~10_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .mask = 16'h048C;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .mask = 16'hECA0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|comb~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .mask = 16'h2E22;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .coord_y = 17;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .mask = 16'h8B0F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Equal3~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .mask = 16'hAAFC;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .mask = 16'h3032;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .mask = 16'h0400;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .mask = 16'h0302;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .mask = 16'h2664;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .mask = 16'hCAC8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .mask = 16'hDDE6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .mask = 16'hFCFE;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(vcc),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .mask = 16'hAA00;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 (
	.A(vcc),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .mask = 16'h000F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~9_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~7_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .mask = 16'hFFF8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~11_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .mask = 16'h5303;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~11_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~12_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .mask = 16'h9810;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~13_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .mask = 16'hFA44;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~13_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~14_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .mask = 16'hDA8A;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|comb~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~15_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .mask = 16'hA280;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~16_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .mask = 16'h88A0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~17_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .mask = 16'h3210;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~15_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~16_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~17_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~18_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .mask = 16'hDDDC;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~18_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~14_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~19_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .mask = 16'h7340;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .mask = 16'h0104;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~20_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .mask = 16'h0A2F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~20_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~19_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~21_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .mask = 16'hCEC2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~22_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .mask = 16'h5410;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~23_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .mask = 16'hA280;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~24_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .mask = 16'h0FAA;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~24_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~25_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .mask = 16'hCCAD;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~26_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .mask = 16'hEE50;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~26_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~27_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .mask = 16'hDAD0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~27_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~25_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~31_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~28_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .mask = 16'hBCB0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~12_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~28_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~21_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~29_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .mask = 16'hF388;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .mask = 16'hECFF;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~23_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~22_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~30_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .mask = 16'h3330;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~30_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~31_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .mask = 16'hC0D1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~3_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .mask = 16'hF020;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .mask = 16'hB020;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .mask = 16'h4F0F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~5_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .mask = 16'hAAA0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .mask = 16'hFC02;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~8_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|comb~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .mask = 16'h32AA;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~5_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~7_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~6_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .mask = 16'h084C;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .mask = 16'hEEFE;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|END~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .mask = 16'h3233;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .mask = 16'h3337;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~2_combout ),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .mask = 16'h000A;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .mask = 16'h4F0F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~4_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~3_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .mask = 16'hFFEC;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SDO~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .mask = 16'h8888;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SDO~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .mask = 16'hFC37;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Equal3~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SDO~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SDO~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .mask = 16'h0501;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Equal5~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SDO~2_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SDO~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .coord_x = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .mask = 16'hCCDC;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|comb~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SDO~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SDO~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .mask = 16'hFD00;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X14_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X14_Y17_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X14_Y17_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y17_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0]~6_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0]~7 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .mask = 16'h55AA;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0]~7 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X14_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X14_Y17_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X14_Y17_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y17_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1]~8_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1]~9 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1]~9 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X14_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X14_Y17_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X14_Y17_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y17_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2]~10_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2]~11 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .mask = 16'hA50A;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2]~11 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X14_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X14_Y17_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X14_Y17_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y17_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3]~13_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3]~14 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3]~14 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X14_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X14_Y17_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X14_Y17_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y17_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4]~15_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4]~16 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4]~16 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X14_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X14_Y17_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X14_Y17_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y17_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~17_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .mask = 16'h3C3C;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SDO~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .mask = 16'h70F0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector2~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .mask = 16'hBFEF;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .mask = 16'h8000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|END~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .mask = 16'hFF13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .mask = 16'h0203;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .mask = 16'h11BB;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~3_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .mask = 16'hF03A;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .mask = 16'h2980;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~5_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .mask = 16'h3939;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .mask = 16'hF858;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector8~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .mask = 16'hBFFB;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector9~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .mask = 16'hFFBE;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(vcc),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Selector9~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector9~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .mask = 16'hFFAA;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|comb~0 (
	.A(vcc),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|comb~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .mask = 16'h00F0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|comb~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|comb~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .coord_y = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .mask = 16'hFD9B;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .mask = 16'h9900;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .mask = 16'h6432;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .mask = 16'hA8A8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .mask = 16'h565A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .mask = 16'h3000;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .mask = 16'h20A0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .mask = 16'hF402;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .mask = 16'h10D0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .mask = 16'hDDD8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .mask = 16'hAB6D;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .mask = 16'hBB0C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .mask = 16'hBBC0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .mask = 16'h5140;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .mask = 16'h30CF;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .mask = 16'hBF88;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .mask = 16'hD000;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .mask = 16'h93B6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .mask = 16'h6BE4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .mask = 16'hDFFE;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .mask = 16'hAF11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .mask = 16'h9D58;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .mask = 16'h0992;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .mask = 16'h936C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .mask = 16'hDDA0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .mask = 16'h5140;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .mask = 16'hEF08;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .mask = 16'hCCED;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .mask = 16'h8A80;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .mask = 16'hC43A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .mask = 16'h4AC8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .mask = 16'h654C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .mask = 16'hA8AD;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .mask = 16'h0082;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .mask = 16'hEE08;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .mask = 16'hD92C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .mask = 16'h6680;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .mask = 16'h53D4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .mask = 16'h3368;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .mask = 16'h5FFE;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .mask = 16'hAB89;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .mask = 16'hD9E0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .mask = 16'hF344;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .mask = 16'h5404;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .mask = 16'hE526;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .mask = 16'h9482;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .mask = 16'h5628;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .mask = 16'h5410;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .mask = 16'h0310;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .mask = 16'hFA44;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .mask = 16'h3D18;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .mask = 16'h5F88;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .mask = 16'h8E3C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .mask = 16'h0801;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .mask = 16'h9102;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .mask = 16'hFF80;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .mask = 16'hB3F6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .mask = 16'h2E10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .mask = 16'hE7F8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .mask = 16'h8CBC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .mask = 16'h1030;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .mask = 16'h7F7C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .mask = 16'h5101;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .mask = 16'hEFBE;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .mask = 16'hFF02;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .mask = 16'hBA98;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .mask = 16'h75BC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .mask = 16'hC7EC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .mask = 16'hFFAE;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .mask = 16'h2406;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .mask = 16'hF50C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .mask = 16'h8226;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .mask = 16'h35F0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .mask = 16'hF838;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .mask = 16'hC8CB;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .mask = 16'h66D4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .coord_x = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .mask = 16'h707A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .mask = 16'hEEEA;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .mask = 16'h0248;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .mask = 16'h001E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .mask = 16'hADA8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .mask = 16'hDCCC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .mask = 16'h0080;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(vcc),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .mask = 16'h5500;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .mask = 16'hD550;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .mask = 16'h51F8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .mask = 16'h0E0C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .mask = 16'hB53F;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .mask = 16'hEDEC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .mask = 16'h3120;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .mask = 16'h231C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .mask = 16'hF303;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .mask = 16'hF3A0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .mask = 16'hB310;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .mask = 16'h92B0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .mask = 16'h98A8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .mask = 16'h5D22;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .mask = 16'h7A70;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .mask = 16'h0B02;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .mask = 16'hF1FE;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .mask = 16'h7B22;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .mask = 16'hA3F0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .mask = 16'h0E02;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .coord_y = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .mask = 16'h2FF6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .mask = 16'hAAD8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .mask = 16'h0708;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .mask = 16'h77C0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .mask = 16'h8CE2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .mask = 16'h2280;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .mask = 16'h3364;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .mask = 16'hF0A3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .mask = 16'hFCFA;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .mask = 16'hFDBC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .mask = 16'h3120;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .mask = 16'hCD89;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .mask = 16'hA680;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .mask = 16'hC460;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .mask = 16'hF6DC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .mask = 16'hE0E5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .mask = 16'h61C8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .mask = 16'h3F88;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .mask = 16'hFF2A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .mask = 16'h182E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .mask = 16'hAAFC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .mask = 16'hC03F;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .mask = 16'h3A88;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .mask = 16'hD3D0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .mask = 16'hF7F0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .coord_x = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .mask = 16'h5F22;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .mask = 16'h68EC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .mask = 16'h7F00;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .mask = 16'hE382;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .coord_x = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .mask = 16'h7B6E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .mask = 16'h6CEC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .mask = 16'hB2EC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .mask = 16'h52F2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .mask = 16'h1032;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .mask = 16'hAEBA;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .mask = 16'hFF10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .mask = 16'h0A70;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .mask = 16'hC03C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .mask = 16'hB834;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .mask = 16'hCBC8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .coord_y = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .mask = 16'hA57E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .mask = 16'h0CC8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .mask = 16'h204C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .mask = 16'h113A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .mask = 16'hCDC1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .mask = 16'h0300;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .mask = 16'h707C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .mask = 16'h1EFC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .mask = 16'hDD2C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .mask = 16'h3FCA;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .coord_y = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .mask = 16'hA800;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .mask = 16'h3090;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .mask = 16'h10E0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .mask = 16'h5804;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .mask = 16'hD020;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .mask = 16'hFE3E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .mask = 16'h46BA;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .mask = 16'hA4AE;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .mask = 16'h0104;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .coord_x = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .coord_y = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .mask = 16'hCAF0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .mask = 16'hB466;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .mask = 16'h2080;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .mask = 16'h006A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .mask = 16'hF0F8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .mask = 16'hE77E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .mask = 16'hB844;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .mask = 16'hFB36;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .mask = 16'hAB89;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .mask = 16'h960A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .coord_x = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .coord_y = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .mask = 16'h53F0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|v_cnt[0] (
	.A(\camera_if_inst|v_cnt [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|v_cnt [0]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[0]~16_combout ),
	.Cout(\camera_if_inst|v_cnt[0]~17 ),
	.Q(\camera_if_inst|v_cnt [0]));
defparam \camera_if_inst|v_cnt[0] .coord_x = 11;
defparam \camera_if_inst|v_cnt[0] .coord_y = 16;
defparam \camera_if_inst|v_cnt[0] .coord_z = 0;
defparam \camera_if_inst|v_cnt[0] .mask = 16'h55AA;
defparam \camera_if_inst|v_cnt[0] .modeMux = 1'b0;
defparam \camera_if_inst|v_cnt[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[0] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[0] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[10] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [10]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[9]~36 ),
	.Qin(\camera_if_inst|v_cnt [10]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[10]~37_combout ),
	.Cout(\camera_if_inst|v_cnt[10]~38 ),
	.Q(\camera_if_inst|v_cnt [10]));
defparam \camera_if_inst|v_cnt[10] .coord_x = 11;
defparam \camera_if_inst|v_cnt[10] .coord_y = 16;
defparam \camera_if_inst|v_cnt[10] .coord_z = 10;
defparam \camera_if_inst|v_cnt[10] .mask = 16'hC30C;
defparam \camera_if_inst|v_cnt[10] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[10] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[10] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[10] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[10] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[11] (
	.A(\camera_if_inst|v_cnt [11]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[10]~38 ),
	.Qin(\camera_if_inst|v_cnt [11]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[11]~39_combout ),
	.Cout(\camera_if_inst|v_cnt[11]~40 ),
	.Q(\camera_if_inst|v_cnt [11]));
defparam \camera_if_inst|v_cnt[11] .coord_x = 11;
defparam \camera_if_inst|v_cnt[11] .coord_y = 16;
defparam \camera_if_inst|v_cnt[11] .coord_z = 11;
defparam \camera_if_inst|v_cnt[11] .mask = 16'h5A5F;
defparam \camera_if_inst|v_cnt[11] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[11] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[11] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[11] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[11] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[12] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [12]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[11]~40 ),
	.Qin(\camera_if_inst|v_cnt [12]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[12]~41_combout ),
	.Cout(\camera_if_inst|v_cnt[12]~42 ),
	.Q(\camera_if_inst|v_cnt [12]));
defparam \camera_if_inst|v_cnt[12] .coord_x = 11;
defparam \camera_if_inst|v_cnt[12] .coord_y = 16;
defparam \camera_if_inst|v_cnt[12] .coord_z = 12;
defparam \camera_if_inst|v_cnt[12] .mask = 16'hC30C;
defparam \camera_if_inst|v_cnt[12] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[12] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[12] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[12] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[12] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[13] (
	.A(\camera_if_inst|v_cnt [13]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[12]~42 ),
	.Qin(\camera_if_inst|v_cnt [13]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[13]~43_combout ),
	.Cout(\camera_if_inst|v_cnt[13]~44 ),
	.Q(\camera_if_inst|v_cnt [13]));
defparam \camera_if_inst|v_cnt[13] .coord_x = 11;
defparam \camera_if_inst|v_cnt[13] .coord_y = 16;
defparam \camera_if_inst|v_cnt[13] .coord_z = 13;
defparam \camera_if_inst|v_cnt[13] .mask = 16'h5A5F;
defparam \camera_if_inst|v_cnt[13] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[13] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[13] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[13] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[13] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[14] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [14]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[13]~44 ),
	.Qin(\camera_if_inst|v_cnt [14]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[14]~45_combout ),
	.Cout(\camera_if_inst|v_cnt[14]~46 ),
	.Q(\camera_if_inst|v_cnt [14]));
defparam \camera_if_inst|v_cnt[14] .coord_x = 11;
defparam \camera_if_inst|v_cnt[14] .coord_y = 16;
defparam \camera_if_inst|v_cnt[14] .coord_z = 14;
defparam \camera_if_inst|v_cnt[14] .mask = 16'hC30C;
defparam \camera_if_inst|v_cnt[14] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[14] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[14] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[14] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[14] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[15] (
	.A(\camera_if_inst|v_cnt [15]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[14]~46 ),
	.Qin(\camera_if_inst|v_cnt [15]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[15]~47_combout ),
	.Cout(),
	.Q(\camera_if_inst|v_cnt [15]));
defparam \camera_if_inst|v_cnt[15] .coord_x = 11;
defparam \camera_if_inst|v_cnt[15] .coord_y = 16;
defparam \camera_if_inst|v_cnt[15] .coord_z = 15;
defparam \camera_if_inst|v_cnt[15] .mask = 16'h5A5A;
defparam \camera_if_inst|v_cnt[15] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[15] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[15] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[15] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[15] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|v_cnt[1] (
	.A(\camera_if_inst|v_cnt [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[0]~17 ),
	.Qin(\camera_if_inst|v_cnt [1]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[1]~19_combout ),
	.Cout(\camera_if_inst|v_cnt[1]~20 ),
	.Q(\camera_if_inst|v_cnt [1]));
defparam \camera_if_inst|v_cnt[1] .coord_x = 11;
defparam \camera_if_inst|v_cnt[1] .coord_y = 16;
defparam \camera_if_inst|v_cnt[1] .coord_z = 1;
defparam \camera_if_inst|v_cnt[1] .mask = 16'h5A5F;
defparam \camera_if_inst|v_cnt[1] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[1] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[1] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[2] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[1]~20 ),
	.Qin(\camera_if_inst|v_cnt [2]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[2]~21_combout ),
	.Cout(\camera_if_inst|v_cnt[2]~22 ),
	.Q(\camera_if_inst|v_cnt [2]));
defparam \camera_if_inst|v_cnt[2] .coord_x = 11;
defparam \camera_if_inst|v_cnt[2] .coord_y = 16;
defparam \camera_if_inst|v_cnt[2] .coord_z = 2;
defparam \camera_if_inst|v_cnt[2] .mask = 16'hC30C;
defparam \camera_if_inst|v_cnt[2] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[2] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[2] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[3] (
	.A(\camera_if_inst|v_cnt [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[2]~22 ),
	.Qin(\camera_if_inst|v_cnt [3]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[3]~23_combout ),
	.Cout(\camera_if_inst|v_cnt[3]~24 ),
	.Q(\camera_if_inst|v_cnt [3]));
defparam \camera_if_inst|v_cnt[3] .coord_x = 11;
defparam \camera_if_inst|v_cnt[3] .coord_y = 16;
defparam \camera_if_inst|v_cnt[3] .coord_z = 3;
defparam \camera_if_inst|v_cnt[3] .mask = 16'h5A5F;
defparam \camera_if_inst|v_cnt[3] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[3] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[3] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[3] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[4] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[3]~24 ),
	.Qin(\camera_if_inst|v_cnt [4]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[4]~25_combout ),
	.Cout(\camera_if_inst|v_cnt[4]~26 ),
	.Q(\camera_if_inst|v_cnt [4]));
defparam \camera_if_inst|v_cnt[4] .coord_x = 11;
defparam \camera_if_inst|v_cnt[4] .coord_y = 16;
defparam \camera_if_inst|v_cnt[4] .coord_z = 4;
defparam \camera_if_inst|v_cnt[4] .mask = 16'hC30C;
defparam \camera_if_inst|v_cnt[4] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[4] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[4] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[5] (
	.A(\camera_if_inst|v_cnt [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[4]~26 ),
	.Qin(\camera_if_inst|v_cnt [5]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[5]~27_combout ),
	.Cout(\camera_if_inst|v_cnt[5]~28 ),
	.Q(\camera_if_inst|v_cnt [5]));
defparam \camera_if_inst|v_cnt[5] .coord_x = 11;
defparam \camera_if_inst|v_cnt[5] .coord_y = 16;
defparam \camera_if_inst|v_cnt[5] .coord_z = 5;
defparam \camera_if_inst|v_cnt[5] .mask = 16'h5A5F;
defparam \camera_if_inst|v_cnt[5] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[5] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[5] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[5] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[6] (
	.A(\camera_if_inst|v_cnt [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[5]~28 ),
	.Qin(\camera_if_inst|v_cnt [6]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[6]~29_combout ),
	.Cout(\camera_if_inst|v_cnt[6]~30 ),
	.Q(\camera_if_inst|v_cnt [6]));
defparam \camera_if_inst|v_cnt[6] .coord_x = 11;
defparam \camera_if_inst|v_cnt[6] .coord_y = 16;
defparam \camera_if_inst|v_cnt[6] .coord_z = 6;
defparam \camera_if_inst|v_cnt[6] .mask = 16'hA50A;
defparam \camera_if_inst|v_cnt[6] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[6] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[6] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[6] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[6] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[7] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[6]~30 ),
	.Qin(\camera_if_inst|v_cnt [7]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[7]~31_combout ),
	.Cout(\camera_if_inst|v_cnt[7]~32 ),
	.Q(\camera_if_inst|v_cnt [7]));
defparam \camera_if_inst|v_cnt[7] .coord_x = 11;
defparam \camera_if_inst|v_cnt[7] .coord_y = 16;
defparam \camera_if_inst|v_cnt[7] .coord_z = 7;
defparam \camera_if_inst|v_cnt[7] .mask = 16'h3C3F;
defparam \camera_if_inst|v_cnt[7] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[7] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[7] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[7] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[7] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[8] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [8]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[7]~32 ),
	.Qin(\camera_if_inst|v_cnt [8]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[8]~33_combout ),
	.Cout(\camera_if_inst|v_cnt[8]~34 ),
	.Q(\camera_if_inst|v_cnt [8]));
defparam \camera_if_inst|v_cnt[8] .coord_x = 11;
defparam \camera_if_inst|v_cnt[8] .coord_y = 16;
defparam \camera_if_inst|v_cnt[8] .coord_z = 8;
defparam \camera_if_inst|v_cnt[8] .mask = 16'hC30C;
defparam \camera_if_inst|v_cnt[8] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[8] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[8] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[8] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[8] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[8]~18 (
	.A(\camera_if_inst|cam_vsync_r [0]),
	.B(\camera_if_inst|Equal3~3_combout ),
	.C(\camera_if_inst|Equal3~2_combout ),
	.D(\camera_if_inst|Equal3~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|v_cnt[8]~18_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|v_cnt[8]~18 .coord_x = 8;
defparam \camera_if_inst|v_cnt[8]~18 .coord_y = 12;
defparam \camera_if_inst|v_cnt[8]~18 .coord_z = 6;
defparam \camera_if_inst|v_cnt[8]~18 .mask = 16'hAAAB;
defparam \camera_if_inst|v_cnt[8]~18 .modeMux = 1'b0;
defparam \camera_if_inst|v_cnt[8]~18 .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[8]~18 .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[8]~18 .BypassEn = 1'b0;
defparam \camera_if_inst|v_cnt[8]~18 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|v_cnt[9] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [9]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[8]~34 ),
	.Qin(\camera_if_inst|v_cnt [9]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X1_Y17_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y17_GND),
	.LutOut(\camera_if_inst|v_cnt[9]~35_combout ),
	.Cout(\camera_if_inst|v_cnt[9]~36 ),
	.Q(\camera_if_inst|v_cnt [9]));
defparam \camera_if_inst|v_cnt[9] .coord_x = 11;
defparam \camera_if_inst|v_cnt[9] .coord_y = 16;
defparam \camera_if_inst|v_cnt[9] .coord_z = 9;
defparam \camera_if_inst|v_cnt[9] .mask = 16'h3C3F;
defparam \camera_if_inst|v_cnt[9] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[9] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[9] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[9] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[9] .CarryEnb = 1'b0;

alta_slice clk_25m(
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\clk_25m~q ),
	.Clk(\e_rxclk~input_o_X33_Y15_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\clk_25m~0_combout ),
	.Cout(),
	.Q(\clk_25m~q ));
defparam clk_25m.coord_x = 46;
defparam clk_25m.coord_y = 15;
defparam clk_25m.coord_z = 15;
defparam clk_25m.mask = 16'h0F0F;
defparam clk_25m.modeMux = 1'b0;
defparam clk_25m.FeedbackMux = 1'b1;
defparam clk_25m.ShiftMux = 1'b0;
defparam clk_25m.BypassEn = 1'b0;
defparam clk_25m.CarryEnb = 1'b1;

alta_io_gclk \clk_25m~clkctrl (
	.inclk(\clk_25m~q ),
	.outclk(\clk_25m~clkctrl_outclk ));
defparam \clk_25m~clkctrl .coord_x = 49;
defparam \clk_25m~clkctrl .coord_y = 15;
defparam \clk_25m~clkctrl .coord_z = 4;

alta_clkenctrl clken_ctrl_X11_Y15_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X11_Y15_SIG_VCC ));
defparam clken_ctrl_X11_Y15_N0.coord_x = 1;
defparam clken_ctrl_X11_Y15_N0.coord_y = 9;
defparam clken_ctrl_X11_Y15_N0.coord_z = 0;
defparam clken_ctrl_X11_Y15_N0.ClkMux = 2'b10;
defparam clken_ctrl_X11_Y15_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X12_Y12_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(reset_init[5]),
	.ClkOut(\clk~inputclkctrl_outclk__reset_init[5]_X12_Y12_SIG_INV ));
defparam clken_ctrl_X12_Y12_N0.coord_x = 47;
defparam clken_ctrl_X12_Y12_N0.coord_y = 15;
defparam clken_ctrl_X12_Y12_N0.coord_z = 0;
defparam clken_ctrl_X12_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X12_Y12_N0.ClkEnMux = 2'b11;

alta_clkenctrl clken_ctrl_X12_Y12_N1(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X12_Y12_SIG_VCC ));
defparam clken_ctrl_X12_Y12_N1.coord_x = 47;
defparam clken_ctrl_X12_Y12_N1.coord_y = 15;
defparam clken_ctrl_X12_Y12_N1.coord_z = 1;
defparam clken_ctrl_X12_Y12_N1.ClkMux = 2'b10;
defparam clken_ctrl_X12_Y12_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X12_Y13_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X12_Y13_SIG_VCC ));
defparam clken_ctrl_X12_Y13_N0.coord_x = 16;
defparam clken_ctrl_X12_Y13_N0.coord_y = 13;
defparam clken_ctrl_X12_Y13_N0.coord_z = 0;
defparam clken_ctrl_X12_Y13_N0.ClkMux = 2'b10;
defparam clken_ctrl_X12_Y13_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X12_Y13_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X12_Y13_SIG_VCC ));
defparam clken_ctrl_X12_Y13_N1.coord_x = 16;
defparam clken_ctrl_X12_Y13_N1.coord_y = 13;
defparam clken_ctrl_X12_Y13_N1.coord_z = 1;
defparam clken_ctrl_X12_Y13_N1.ClkMux = 2'b10;
defparam clken_ctrl_X12_Y13_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X12_Y14_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ));
defparam clken_ctrl_X12_Y14_N0.coord_x = 2;
defparam clken_ctrl_X12_Y14_N0.coord_y = 9;
defparam clken_ctrl_X12_Y14_N0.coord_z = 0;
defparam clken_ctrl_X12_Y14_N0.ClkMux = 2'b10;
defparam clken_ctrl_X12_Y14_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X12_Y15_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ));
defparam clken_ctrl_X12_Y15_N0.coord_x = 2;
defparam clken_ctrl_X12_Y15_N0.coord_y = 10;
defparam clken_ctrl_X12_Y15_N0.coord_z = 0;
defparam clken_ctrl_X12_Y15_N0.ClkMux = 2'b10;
defparam clken_ctrl_X12_Y15_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X13_Y12_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X13_Y12_SIG_VCC ));
defparam clken_ctrl_X13_Y12_N0.coord_x = 15;
defparam clken_ctrl_X13_Y12_N0.coord_y = 16;
defparam clken_ctrl_X13_Y12_N0.coord_z = 0;
defparam clken_ctrl_X13_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X13_Y12_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X13_Y12_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X13_Y12_SIG_VCC ));
defparam clken_ctrl_X13_Y12_N1.coord_x = 15;
defparam clken_ctrl_X13_Y12_N1.coord_y = 16;
defparam clken_ctrl_X13_Y12_N1.coord_z = 1;
defparam clken_ctrl_X13_Y12_N1.ClkMux = 2'b10;
defparam clken_ctrl_X13_Y12_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X13_Y13_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout ),
	.ClkOut(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X13_Y13_SIG_SIG ));
defparam clken_ctrl_X13_Y13_N0.coord_x = 15;
defparam clken_ctrl_X13_Y13_N0.coord_y = 13;
defparam clken_ctrl_X13_Y13_N0.coord_z = 0;
defparam clken_ctrl_X13_Y13_N0.ClkMux = 2'b10;
defparam clken_ctrl_X13_Y13_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X13_Y13_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X13_Y13_SIG_VCC ));
defparam clken_ctrl_X13_Y13_N1.coord_x = 15;
defparam clken_ctrl_X13_Y13_N1.coord_y = 13;
defparam clken_ctrl_X13_Y13_N1.coord_z = 1;
defparam clken_ctrl_X13_Y13_N1.ClkMux = 2'b10;
defparam clken_ctrl_X13_Y13_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X14_Y12_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y12_SIG_SIG ));
defparam clken_ctrl_X14_Y12_N0.coord_x = 17;
defparam clken_ctrl_X14_Y12_N0.coord_y = 16;
defparam clken_ctrl_X14_Y12_N0.coord_z = 0;
defparam clken_ctrl_X14_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y12_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X14_Y12_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X14_Y12_SIG_VCC ));
defparam clken_ctrl_X14_Y12_N1.coord_x = 17;
defparam clken_ctrl_X14_Y12_N1.coord_y = 16;
defparam clken_ctrl_X14_Y12_N1.coord_z = 1;
defparam clken_ctrl_X14_Y12_N1.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y12_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X14_Y13_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ClkOut(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y13_SIG_SIG ));
defparam clken_ctrl_X14_Y13_N0.coord_x = 17;
defparam clken_ctrl_X14_Y13_N0.coord_y = 13;
defparam clken_ctrl_X14_Y13_N0.coord_z = 0;
defparam clken_ctrl_X14_Y13_N0.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y13_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X14_Y13_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X14_Y13_SIG_VCC ));
defparam clken_ctrl_X14_Y13_N1.coord_x = 17;
defparam clken_ctrl_X14_Y13_N1.coord_y = 13;
defparam clken_ctrl_X14_Y13_N1.coord_z = 1;
defparam clken_ctrl_X14_Y13_N1.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y13_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X14_Y17_N1(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X14_Y17_SIG_SIG ));
defparam clken_ctrl_X14_Y17_N1.coord_x = 10;
defparam clken_ctrl_X14_Y17_N1.coord_y = 15;
defparam clken_ctrl_X14_Y17_N1.coord_z = 1;
defparam clken_ctrl_X14_Y17_N1.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y17_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y11_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X16_Y11_SIG_VCC ));
defparam clken_ctrl_X16_Y11_N0.coord_x = 17;
defparam clken_ctrl_X16_Y11_N0.coord_y = 15;
defparam clken_ctrl_X16_Y11_N0.coord_z = 0;
defparam clken_ctrl_X16_Y11_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y11_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X16_Y11_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y11_SIG_SIG ));
defparam clken_ctrl_X16_Y11_N1.coord_x = 17;
defparam clken_ctrl_X16_Y11_N1.coord_y = 15;
defparam clken_ctrl_X16_Y11_N1.coord_z = 1;
defparam clken_ctrl_X16_Y11_N1.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y11_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y12_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ));
defparam clken_ctrl_X16_Y12_N0.coord_x = 16;
defparam clken_ctrl_X16_Y12_N0.coord_y = 16;
defparam clken_ctrl_X16_Y12_N0.coord_z = 0;
defparam clken_ctrl_X16_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y12_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X16_Y12_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y12_SIG_SIG ));
defparam clken_ctrl_X16_Y12_N1.coord_x = 16;
defparam clken_ctrl_X16_Y12_N1.coord_y = 16;
defparam clken_ctrl_X16_Y12_N1.coord_z = 1;
defparam clken_ctrl_X16_Y12_N1.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y12_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y13_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ClkOut(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y13_SIG_SIG ));
defparam clken_ctrl_X16_Y13_N0.coord_x = 17;
defparam clken_ctrl_X16_Y13_N0.coord_y = 14;
defparam clken_ctrl_X16_Y13_N0.coord_z = 0;
defparam clken_ctrl_X16_Y13_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y13_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y13_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X16_Y13_SIG_VCC ));
defparam clken_ctrl_X16_Y13_N1.coord_x = 17;
defparam clken_ctrl_X16_Y13_N1.coord_y = 14;
defparam clken_ctrl_X16_Y13_N1.coord_z = 1;
defparam clken_ctrl_X16_Y13_N1.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y13_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X16_Y16_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y16_SIG_SIG ));
defparam clken_ctrl_X16_Y16_N0.coord_x = 11;
defparam clken_ctrl_X16_Y16_N0.coord_y = 15;
defparam clken_ctrl_X16_Y16_N0.coord_z = 0;
defparam clken_ctrl_X16_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y16_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y17_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y17_SIG_SIG ));
defparam clken_ctrl_X16_Y17_N0.coord_x = 10;
defparam clken_ctrl_X16_Y17_N0.coord_y = 13;
defparam clken_ctrl_X16_Y17_N0.coord_z = 0;
defparam clken_ctrl_X16_Y17_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y17_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y18_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y18_SIG_SIG ));
defparam clken_ctrl_X16_Y18_N0.coord_x = 11;
defparam clken_ctrl_X16_Y18_N0.coord_y = 14;
defparam clken_ctrl_X16_Y18_N0.coord_z = 0;
defparam clken_ctrl_X16_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y18_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X17_Y12_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X17_Y12_SIG_VCC ));
defparam clken_ctrl_X17_Y12_N0.coord_x = 15;
defparam clken_ctrl_X17_Y12_N0.coord_y = 15;
defparam clken_ctrl_X17_Y12_N0.coord_z = 0;
defparam clken_ctrl_X17_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y12_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y13_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X17_Y13_SIG_VCC ));
defparam clken_ctrl_X17_Y13_N0.coord_x = 16;
defparam clken_ctrl_X17_Y13_N0.coord_y = 15;
defparam clken_ctrl_X17_Y13_N0.coord_z = 0;
defparam clken_ctrl_X17_Y13_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y13_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y13_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X17_Y13_SIG_VCC ));
defparam clken_ctrl_X17_Y13_N1.coord_x = 16;
defparam clken_ctrl_X17_Y13_N1.coord_y = 15;
defparam clken_ctrl_X17_Y13_N1.coord_z = 1;
defparam clken_ctrl_X17_Y13_N1.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y13_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y14_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X17_Y14_SIG_VCC ));
defparam clken_ctrl_X17_Y14_N0.coord_x = 16;
defparam clken_ctrl_X17_Y14_N0.coord_y = 14;
defparam clken_ctrl_X17_Y14_N0.coord_z = 0;
defparam clken_ctrl_X17_Y14_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y14_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y17_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y17_SIG_SIG ));
defparam clken_ctrl_X17_Y17_N0.coord_x = 11;
defparam clken_ctrl_X17_Y17_N0.coord_y = 13;
defparam clken_ctrl_X17_Y17_N0.coord_z = 0;
defparam clken_ctrl_X17_Y17_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y17_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X17_Y17_N1(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X17_Y17_SIG_VCC ));
defparam clken_ctrl_X17_Y17_N1.coord_x = 11;
defparam clken_ctrl_X17_Y17_N1.coord_y = 13;
defparam clken_ctrl_X17_Y17_N1.coord_z = 1;
defparam clken_ctrl_X17_Y17_N1.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y17_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y1_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked ),
	.ClkEn(),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked_X17_Y1_SIG_VCC ));
defparam clken_ctrl_X17_Y1_N0.coord_x = 1;
defparam clken_ctrl_X17_Y1_N0.coord_y = 1;
defparam clken_ctrl_X17_Y1_N0.coord_z = 0;
defparam clken_ctrl_X17_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y1_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X18_Y17_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y17_SIG_SIG ));
defparam clken_ctrl_X18_Y17_N0.coord_x = 13;
defparam clken_ctrl_X18_Y17_N0.coord_y = 13;
defparam clken_ctrl_X18_Y17_N0.coord_z = 0;
defparam clken_ctrl_X18_Y17_N0.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y17_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X18_Y17_N1(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X18_Y17_SIG_SIG ));
defparam clken_ctrl_X18_Y17_N1.coord_x = 13;
defparam clken_ctrl_X18_Y17_N1.coord_y = 13;
defparam clken_ctrl_X18_Y17_N1.coord_z = 1;
defparam clken_ctrl_X18_Y17_N1.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y17_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X19_Y12_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout_X19_Y12_SIG_SIG ));
defparam clken_ctrl_X19_Y12_N0.coord_x = 19;
defparam clken_ctrl_X19_Y12_N0.coord_y = 16;
defparam clken_ctrl_X19_Y12_N0.coord_z = 0;
defparam clken_ctrl_X19_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X19_Y12_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X1_Y17_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(\camera_if_inst|v_cnt[8]~18_combout ),
	.ClkOut(\cam_pclk~input_o__camera_if_inst|v_cnt[8]~18_combout_X1_Y17_SIG_SIG ));
defparam clken_ctrl_X1_Y17_N1.coord_x = 11;
defparam clken_ctrl_X1_Y17_N1.coord_y = 16;
defparam clken_ctrl_X1_Y17_N1.coord_z = 1;
defparam clken_ctrl_X1_Y17_N1.ClkMux = 2'b10;
defparam clken_ctrl_X1_Y17_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X1_Y7_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X1_Y7_SIG_VCC ));
defparam clken_ctrl_X1_Y7_N0.coord_x = 8;
defparam clken_ctrl_X1_Y7_N0.coord_y = 12;
defparam clken_ctrl_X1_Y7_N0.coord_z = 0;
defparam clken_ctrl_X1_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X1_Y7_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X21_Y18_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|crc32_inst|crc_data[28]~9_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ));
defparam clken_ctrl_X21_Y18_N0.coord_x = 20;
defparam clken_ctrl_X21_Y18_N0.coord_y = 16;
defparam clken_ctrl_X21_Y18_N0.coord_z = 0;
defparam clken_ctrl_X21_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X21_Y18_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X21_Y19_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|crc32_inst|crc_data[28]~9_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y19_SIG_SIG ));
defparam clken_ctrl_X21_Y19_N0.coord_x = 20;
defparam clken_ctrl_X21_Y19_N0.coord_y = 17;
defparam clken_ctrl_X21_Y19_N0.coord_z = 0;
defparam clken_ctrl_X21_Y19_N0.ClkMux = 2'b10;
defparam clken_ctrl_X21_Y19_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X22_Y16_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X22_Y16_SIG_SIG ));
defparam clken_ctrl_X22_Y16_N1.coord_x = 22;
defparam clken_ctrl_X22_Y16_N1.coord_y = 16;
defparam clken_ctrl_X22_Y16_N1.coord_z = 1;
defparam clken_ctrl_X22_Y16_N1.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y16_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X22_Y19_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|crc32_inst|crc_data[28]~9_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X22_Y19_SIG_SIG ));
defparam clken_ctrl_X22_Y19_N0.coord_x = 19;
defparam clken_ctrl_X22_Y19_N0.coord_y = 17;
defparam clken_ctrl_X22_Y19_N0.coord_z = 0;
defparam clken_ctrl_X22_Y19_N0.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y19_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X22_Y19_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X22_Y19_SIG_VCC ));
defparam clken_ctrl_X22_Y19_N1.coord_x = 19;
defparam clken_ctrl_X22_Y19_N1.coord_y = 17;
defparam clken_ctrl_X22_Y19_N1.coord_z = 1;
defparam clken_ctrl_X22_Y19_N1.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y19_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X22_Y8_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X22_Y8_SIG_VCC ));
defparam clken_ctrl_X22_Y8_N0.coord_x = 10;
defparam clken_ctrl_X22_Y8_N0.coord_y = 17;
defparam clken_ctrl_X22_Y8_N0.coord_z = 0;
defparam clken_ctrl_X22_Y8_N0.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y8_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X23_Y15_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ));
defparam clken_ctrl_X23_Y15_N1.coord_x = 22;
defparam clken_ctrl_X23_Y15_N1.coord_y = 18;
defparam clken_ctrl_X23_Y15_N1.coord_z = 1;
defparam clken_ctrl_X23_Y15_N1.ClkMux = 2'b10;
defparam clken_ctrl_X23_Y15_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X23_Y16_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X23_Y16_SIG_VCC ));
defparam clken_ctrl_X23_Y16_N0.coord_x = 21;
defparam clken_ctrl_X23_Y16_N0.coord_y = 13;
defparam clken_ctrl_X23_Y16_N0.coord_z = 0;
defparam clken_ctrl_X23_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X23_Y16_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X23_Y16_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y16_SIG_SIG ));
defparam clken_ctrl_X23_Y16_N1.coord_x = 21;
defparam clken_ctrl_X23_Y16_N1.coord_y = 13;
defparam clken_ctrl_X23_Y16_N1.coord_z = 1;
defparam clken_ctrl_X23_Y16_N1.ClkMux = 2'b10;
defparam clken_ctrl_X23_Y16_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X23_Y18_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X23_Y18_SIG_VCC ));
defparam clken_ctrl_X23_Y18_N0.coord_x = 21;
defparam clken_ctrl_X23_Y18_N0.coord_y = 16;
defparam clken_ctrl_X23_Y18_N0.coord_z = 0;
defparam clken_ctrl_X23_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X23_Y18_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X23_Y18_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y18_SIG_SIG ));
defparam clken_ctrl_X23_Y18_N1.coord_x = 21;
defparam clken_ctrl_X23_Y18_N1.coord_y = 16;
defparam clken_ctrl_X23_Y18_N1.coord_z = 1;
defparam clken_ctrl_X23_Y18_N1.ClkMux = 2'b10;
defparam clken_ctrl_X23_Y18_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X23_Y19_N0(
	.ClkIn(\e_rxclk~input_o ),
	.ClkEn(),
	.ClkOut(\e_rxclk~input_o_X23_Y19_INV_VCC ));
defparam clken_ctrl_X23_Y19_N0.coord_x = 21;
defparam clken_ctrl_X23_Y19_N0.coord_y = 17;
defparam clken_ctrl_X23_Y19_N0.coord_z = 0;
defparam clken_ctrl_X23_Y19_N0.ClkMux = 2'b11;
defparam clken_ctrl_X23_Y19_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X23_Y19_N1(
	.ClkIn(\e_rxclk~input_o ),
	.ClkEn(\mii_to_rmii_inst|tx_dv_reg~q ),
	.ClkOut(\e_rxclk~input_o__mii_to_rmii_inst|tx_dv_reg~q_X23_Y19_SIG_SIG ));
defparam clken_ctrl_X23_Y19_N1.coord_x = 21;
defparam clken_ctrl_X23_Y19_N1.coord_y = 17;
defparam clken_ctrl_X23_Y19_N1.coord_z = 1;
defparam clken_ctrl_X23_Y19_N1.ClkMux = 2'b10;
defparam clken_ctrl_X23_Y19_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X23_Y8_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X23_Y8_SIG_VCC ));
defparam clken_ctrl_X23_Y8_N0.coord_x = 11;
defparam clken_ctrl_X23_Y8_N0.coord_y = 17;
defparam clken_ctrl_X23_Y8_N0.coord_z = 0;
defparam clken_ctrl_X23_Y8_N0.ClkMux = 2'b10;
defparam clken_ctrl_X23_Y8_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X24_Y15_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X24_Y15_SIG_VCC ));
defparam clken_ctrl_X24_Y15_N0.coord_x = 20;
defparam clken_ctrl_X24_Y15_N0.coord_y = 15;
defparam clken_ctrl_X24_Y15_N0.coord_z = 0;
defparam clken_ctrl_X24_Y15_N0.ClkMux = 2'b10;
defparam clken_ctrl_X24_Y15_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X24_Y15_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X24_Y15_SIG_SIG ));
defparam clken_ctrl_X24_Y15_N1.coord_x = 20;
defparam clken_ctrl_X24_Y15_N1.coord_y = 15;
defparam clken_ctrl_X24_Y15_N1.coord_z = 1;
defparam clken_ctrl_X24_Y15_N1.ClkMux = 2'b10;
defparam clken_ctrl_X24_Y15_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X24_Y16_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|cnt[3]~13_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[3]~13_combout_X24_Y16_SIG_SIG ));
defparam clken_ctrl_X24_Y16_N1.coord_x = 22;
defparam clken_ctrl_X24_Y16_N1.coord_y = 14;
defparam clken_ctrl_X24_Y16_N1.coord_z = 1;
defparam clken_ctrl_X24_Y16_N1.ClkMux = 2'b10;
defparam clken_ctrl_X24_Y16_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X25_Y16_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X25_Y16_SIG_SIG ));
defparam clken_ctrl_X25_Y16_N0.coord_x = 21;
defparam clken_ctrl_X25_Y16_N0.coord_y = 14;
defparam clken_ctrl_X25_Y16_N0.coord_z = 0;
defparam clken_ctrl_X25_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X25_Y16_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X25_Y16_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X25_Y16_SIG_VCC ));
defparam clken_ctrl_X25_Y16_N1.coord_x = 21;
defparam clken_ctrl_X25_Y16_N1.coord_y = 14;
defparam clken_ctrl_X25_Y16_N1.coord_z = 1;
defparam clken_ctrl_X25_Y16_N1.ClkMux = 2'b10;
defparam clken_ctrl_X25_Y16_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X25_Y17_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|always3~4_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ));
defparam clken_ctrl_X25_Y17_N0.coord_x = 19;
defparam clken_ctrl_X25_Y17_N0.coord_y = 11;
defparam clken_ctrl_X25_Y17_N0.coord_z = 0;
defparam clken_ctrl_X25_Y17_N0.ClkMux = 2'b10;
defparam clken_ctrl_X25_Y17_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X28_Y14_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|check_sum[8]~47_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y14_SIG_SIG ));
defparam clken_ctrl_X28_Y14_N0.coord_x = 21;
defparam clken_ctrl_X28_Y14_N0.coord_y = 9;
defparam clken_ctrl_X28_Y14_N0.coord_z = 0;
defparam clken_ctrl_X28_Y14_N0.ClkMux = 2'b10;
defparam clken_ctrl_X28_Y14_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X28_Y14_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y14_SIG_SIG ));
defparam clken_ctrl_X28_Y14_N1.coord_x = 21;
defparam clken_ctrl_X28_Y14_N1.coord_y = 9;
defparam clken_ctrl_X28_Y14_N1.coord_z = 1;
defparam clken_ctrl_X28_Y14_N1.ClkMux = 2'b10;
defparam clken_ctrl_X28_Y14_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X28_Y15_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y15_SIG_SIG ));
defparam clken_ctrl_X28_Y15_N0.coord_x = 21;
defparam clken_ctrl_X28_Y15_N0.coord_y = 10;
defparam clken_ctrl_X28_Y15_N0.coord_z = 0;
defparam clken_ctrl_X28_Y15_N0.ClkMux = 2'b10;
defparam clken_ctrl_X28_Y15_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X28_Y15_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|check_sum[8]~47_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y15_SIG_SIG ));
defparam clken_ctrl_X28_Y15_N1.coord_x = 21;
defparam clken_ctrl_X28_Y15_N1.coord_y = 10;
defparam clken_ctrl_X28_Y15_N1.coord_z = 1;
defparam clken_ctrl_X28_Y15_N1.ClkMux = 2'b10;
defparam clken_ctrl_X28_Y15_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X28_Y18_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y18_SIG_SIG ));
defparam clken_ctrl_X28_Y18_N0.coord_x = 20;
defparam clken_ctrl_X28_Y18_N0.coord_y = 10;
defparam clken_ctrl_X28_Y18_N0.coord_z = 0;
defparam clken_ctrl_X28_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X28_Y18_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X2_Y7_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X2_Y7_SIG_VCC ));
defparam clken_ctrl_X2_Y7_N0.coord_x = 9;
defparam clken_ctrl_X2_Y7_N0.coord_y = 12;
defparam clken_ctrl_X2_Y7_N0.coord_z = 0;
defparam clken_ctrl_X2_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X2_Y7_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X33_Y15_N0(
	.ClkIn(\e_rxclk~input_o ),
	.ClkEn(),
	.ClkOut(\e_rxclk~input_o_X33_Y15_INV_VCC ));
defparam clken_ctrl_X33_Y15_N0.coord_x = 46;
defparam clken_ctrl_X33_Y15_N0.coord_y = 15;
defparam clken_ctrl_X33_Y15_N0.coord_z = 0;
defparam clken_ctrl_X33_Y15_N0.ClkMux = 2'b11;
defparam clken_ctrl_X33_Y15_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X3_Y7_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X3_Y7_SIG_VCC ));
defparam clken_ctrl_X3_Y7_N0.coord_x = 14;
defparam clken_ctrl_X3_Y7_N0.coord_y = 16;
defparam clken_ctrl_X3_Y7_N0.coord_z = 0;
defparam clken_ctrl_X3_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X3_Y7_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X3_Y7_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X3_Y7_SIG_VCC ));
defparam clken_ctrl_X3_Y7_N1.coord_x = 14;
defparam clken_ctrl_X3_Y7_N1.coord_y = 16;
defparam clken_ctrl_X3_Y7_N1.coord_z = 1;
defparam clken_ctrl_X3_Y7_N1.ClkMux = 2'b10;
defparam clken_ctrl_X3_Y7_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X4_Y7_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X4_Y7_SIG_VCC ));
defparam clken_ctrl_X4_Y7_N0.coord_x = 17;
defparam clken_ctrl_X4_Y7_N0.coord_y = 12;
defparam clken_ctrl_X4_Y7_N0.coord_z = 0;
defparam clken_ctrl_X4_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X4_Y7_N0.ClkEnMux = 2'b01;

alta_dio \clk~input (
	.padio(clk),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\clk~input_o ),
	.regout());
defparam \clk~input .coord_x = 0;
defparam \clk~input .coord_y = 12;
defparam \clk~input .coord_z = 2;
defparam \clk~input .IN_ASYNC_MODE = 1'b0;
defparam \clk~input .IN_SYNC_MODE = 1'b0;
defparam \clk~input .IN_POWERUP = 1'b0;
defparam \clk~input .IN_ASYNC_DISABLE = 1'b0;
defparam \clk~input .IN_SYNC_DISABLE = 1'b0;
defparam \clk~input .OUT_REG_MODE = 1'b0;
defparam \clk~input .OUT_ASYNC_MODE = 1'b0;
defparam \clk~input .OUT_SYNC_MODE = 1'b0;
defparam \clk~input .OUT_POWERUP = 1'b0;
defparam \clk~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \clk~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \clk~input .OUT_SYNC_DISABLE = 1'b0;
defparam \clk~input .OUT_DDIO = 1'b0;
defparam \clk~input .OE_REG_MODE = 1'b0;
defparam \clk~input .OE_ASYNC_MODE = 1'b0;
defparam \clk~input .OE_SYNC_MODE = 1'b0;
defparam \clk~input .OE_POWERUP = 1'b0;
defparam \clk~input .OE_CLKEN_DISABLE = 1'b0;
defparam \clk~input .OE_ASYNC_DISABLE = 1'b0;
defparam \clk~input .OE_SYNC_DISABLE = 1'b0;
defparam \clk~input .OE_DDIO = 1'b0;
defparam \clk~input .CFG_TRI_INPUT = 1'b0;
defparam \clk~input .CFG_PULL_UP = 1'b0;
defparam \clk~input .CFG_OPEN_DRAIN = 1'b0;
defparam \clk~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \clk~input .CFG_PDRV = 7'b0010000;
defparam \clk~input .CFG_NDRV = 7'b0010000;
defparam \clk~input .CFG_KEEP = 2'b00;
defparam \clk~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \clk~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \clk~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \clk~input .CFG_LVDS_IN_EN = 1'b0;
defparam \clk~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \clk~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \clk~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \clk~input .CFG_OSCDIV = 2'b00;
defparam \clk~input .CFG_ROCTUSR = 1'b0;
defparam \clk~input .CFG_SEL_CUA = 1'b0;
defparam \clk~input .CFG_ROCT_EN = 1'b0;
defparam \clk~input .INPUT_ONLY = 1'b1;
defparam \clk~input .DPCLK_DELAY = 4'b0000;
defparam \clk~input .OUT_DELAY = 1'b0;
defparam \clk~input .IN_DATA_DELAY = 3'b000;
defparam \clk~input .IN_REG_DELAY = 3'b000;

alta_io_gclk \clk~inputclkctrl (
	.inclk(\clk~input_o ),
	.outclk(\clk~inputclkctrl_outclk ));
defparam \clk~inputclkctrl .coord_x = 0;
defparam \clk~inputclkctrl .coord_y = 12;
defparam \clk~inputclkctrl .coord_z = 0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .mask = 16'hF000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~COUT ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .mask = 16'h0F0F;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [0]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita0~combout ),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita0~COUT ),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .mask = 16'h3333;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita0~COUT ),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [1]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~combout ),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~COUT ),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .mask = 16'h5A5F;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [0]),
	.Clk(\cam_pclk~input_o_X3_Y7_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X3_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .coord_x = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [12]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [10]),
	.Clk(\cam_pclk~input_o_X16_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [1]),
	.Clk(\cam_pclk~input_o_X13_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ),
	.SyncReset(SyncReset_X13_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y12_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [2]),
	.Clk(\cam_pclk~input_o_X12_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [3]),
	.Clk(\cam_pclk~input_o_X3_Y7_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X3_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .coord_x = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [4]),
	.Clk(\cam_pclk~input_o_X13_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [5]),
	.Clk(\cam_pclk~input_o_X12_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [6]),
	.Clk(\cam_pclk~input_o_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [7]),
	.Clk(\cam_pclk~input_o_X13_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ),
	.SyncReset(SyncReset_X13_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y12_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [8]),
	.Clk(\cam_pclk~input_o_X16_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(SyncReset_X16_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y13_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [11]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [9]),
	.Clk(\cam_pclk~input_o_X16_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .CarryEnb = 1'b1;

alta_bram9k \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 (
	.DataInA({vcc, \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], vcc, \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0]}),
	.DataInB({1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz}),
	.AddressA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0], vcc}),
	.AddressB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0_combout , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell_combout , vcc, vcc, vcc}),
	.ByteEnA({vcc, vcc}),
	.ByteEnB({1'bz, 1'bz}),
	.DataOutA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [0]}),
	.DataOutB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [0]}),
	.Clk0(\cam_pclk~input_o ),
	.ClkEn0(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.AsyncReset0(gnd),
	.Clk1(\clk_25m~clkctrl_outclk ),
	.ClkEn1(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.AsyncReset1(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.WeA(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ReA(gnd),
	.WeB(gnd),
	.ReB(vcc),
	.AddressStallA(gnd),
	.AddressStallB(!\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .coord_x = 18;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .CLKMODE = 2'b10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PACKEDMODE = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_CLKIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_CLKOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_CLKIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_CLKOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_RSTIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_RSTOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_RSTIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_RSTOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_WIDTH = 5'b01110;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_WIDTH = 5'b01000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_OUTREG = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_OUTREG = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .RSEN_DLY = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .DLYTIME = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .INIT_VAL = 9216'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

alta_bram9k \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 (
	.DataInA({vcc, \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [1], \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [1], \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [1], \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [1], vcc, \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [1], \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [1], \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [1], \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [1]}),
	.DataInB({1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz}),
	.AddressA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0], vcc}),
	.AddressB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0_combout , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell_combout , vcc, vcc, vcc}),
	.ByteEnA({vcc, vcc}),
	.ByteEnB({1'bz, 1'bz}),
	.DataOutA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [0]}),
	.DataOutB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [0]}),
	.Clk0(\cam_pclk~input_o ),
	.ClkEn0(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.AsyncReset0(gnd),
	.Clk1(\clk_25m~clkctrl_outclk ),
	.ClkEn1(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.AsyncReset1(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.WeA(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ReA(gnd),
	.WeB(gnd),
	.ReB(vcc),
	.AddressStallA(gnd),
	.AddressStallB(!\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .coord_x = 18;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .CLKMODE = 2'b10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PACKEDMODE = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_CLKIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_CLKOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_CLKIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_CLKOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_RSTIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_RSTOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_RSTIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_RSTOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_WIDTH = 5'b01110;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_WIDTH = 5'b01000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_OUTREG = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_OUTREG = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .RSEN_DLY = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .DLYTIME = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .INIT_VAL = 9216'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

alta_bram9k \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 (
	.DataInA({vcc, \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [2], \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [2], \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [2], \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [2], vcc, \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [2], \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [2], \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [2], \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [2]}),
	.DataInB({1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz}),
	.AddressA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0], vcc}),
	.AddressB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0_combout , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell_combout , vcc, vcc, vcc}),
	.ByteEnA({vcc, vcc}),
	.ByteEnB({1'bz, 1'bz}),
	.DataOutA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [0]}),
	.DataOutB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [0]}),
	.Clk0(\cam_pclk~input_o ),
	.ClkEn0(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.AsyncReset0(gnd),
	.Clk1(\clk_25m~clkctrl_outclk ),
	.ClkEn1(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.AsyncReset1(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.WeA(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ReA(gnd),
	.WeB(gnd),
	.ReB(vcc),
	.AddressStallA(gnd),
	.AddressStallB(!\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .coord_x = 18;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .CLKMODE = 2'b10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PACKEDMODE = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_CLKIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_CLKOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_CLKIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_CLKOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_RSTIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_RSTOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_RSTIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_RSTOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_WIDTH = 5'b01110;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_WIDTH = 5'b01000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_OUTREG = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_OUTREG = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .RSEN_DLY = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .DLYTIME = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .INIT_VAL = 9216'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

alta_bram9k \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 (
	.DataInA({vcc, \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [3], vcc, \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [3]}),
	.DataInB({1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz}),
	.AddressA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0], vcc}),
	.AddressB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0_combout , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell_combout , vcc, vcc, vcc}),
	.ByteEnA({vcc, vcc}),
	.ByteEnB({1'bz, 1'bz}),
	.DataOutA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutA [0]}),
	.DataOutB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [0]}),
	.Clk0(\cam_pclk~input_o ),
	.ClkEn0(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.AsyncReset0(gnd),
	.Clk1(\clk_25m~clkctrl_outclk ),
	.ClkEn1(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.AsyncReset1(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.WeA(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ReA(gnd),
	.WeB(gnd),
	.ReB(vcc),
	.AddressStallA(gnd),
	.AddressStallB(!\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .coord_x = 18;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .CLKMODE = 2'b10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PACKEDMODE = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTA_CLKIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTA_CLKOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTB_CLKIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTB_CLKOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTA_RSTIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTA_RSTOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTB_RSTIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTB_RSTOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTA_WIDTH = 5'b01110;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTB_WIDTH = 5'b01000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTA_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTB_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTA_OUTREG = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .PORTB_OUTREG = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .RSEN_DLY = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .DLYTIME = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3 .INIT_VAL = 9216'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [0]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1_cout ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .mask = 16'h00DD;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [5]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11_cout ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .mask = 16'h004D;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [6]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [6]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12_combout ),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~13 ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .mask = 16'h962B;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [7]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14_combout ),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~15 ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .mask = 16'h694D;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [8]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [8]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16_combout ),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~17 ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .mask = 16'h964D;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [9]),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [9]),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .mask = 16'h5AA5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [1]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3_cout ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .mask = 16'h004D;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [2]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5_cout ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .mask = 16'h002B;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [3]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7_cout ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .mask = 16'h004D;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [4]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9_cout ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .mask = 16'h004D;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~1_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~0_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~3_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .mask = 16'hFFFE;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .mask = 16'h6666;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .mask = 16'h2000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .mask = 16'h1000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .mask = 16'h0400;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .mask = 16'h0200;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .mask = 16'h0004;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .mask = 16'h0100;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y12_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~1_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .mask = 16'h3C3C;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .mask = 16'h00FF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .mask = 16'hF0D2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~q ),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y11_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .mask = 16'hB4B4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .mask = 16'h0FF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .mask = 16'h3CF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .mask = 16'hD2F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .mask = 16'h5A5A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y11_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .mask = 16'h5AF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y11_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .mask = 16'hB4F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y11_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .mask = 16'h0FF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~q ),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y11_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .mask = 16'h7878;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [1]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [0]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [2]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y12_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~7_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .mask = 16'h6699;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [0]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y12_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~10_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .mask = 16'h9669;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [1]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y12_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~9_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [2]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~8_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .mask = 16'h9966;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [0]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y12_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .mask = 16'h00FF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~q ),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(SyncReset_X16_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y11_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [1]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y12_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y12_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y12_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(SyncReset_X16_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y12_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [4]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y12_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y12_SIG ),
	.SyncReset(SyncReset_X14_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y12_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(SyncReset_X16_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y11_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [7]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~q ),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(SyncReset_X16_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y11_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor1~combout ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [0]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [0]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor0~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .mask = 16'h33CC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor4~combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [1]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [1]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor1~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor4~combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [2]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor2~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .mask = 16'h9696;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor4~combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [3]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor3~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .mask = 16'h3C3C;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [4]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor7~combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [4]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor4~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5]),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor7~combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [5]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor5~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .mask = 16'hA55A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor7~combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [6]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor6~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .mask = 16'h0FF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [7]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [7]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor7~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8]),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [8]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor8~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .mask = 16'hA55A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [9]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y11_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor9~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .mask = 16'h6666;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [0]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor1~combout ),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [0]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor0~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .mask = 16'h3C3C;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [2]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [1]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor4~combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [1]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor1~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [2]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor4~combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [2]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor2~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .mask = 16'hC33C;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor4~combout ),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [3]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor3~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .mask = 16'h55AA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [4]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [5]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor7~combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [6]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [4]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor4~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [6]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor7~combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [5]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [5]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor5~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .mask = 16'hC33C;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor7~combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [6]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [6]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor6~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .mask = 16'h0FF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [7]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [8]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [7]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor7~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [8]),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [8]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor8~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .mask = 16'hA55A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [9]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor9~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .mask = 16'h3C3C;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [0]),
	.Clk(\clk_25m~clkctrl_outclk_X3_Y7_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X3_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .coord_x = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [10]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [10]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y14_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [1]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [1]),
	.Clk(\clk_25m~clkctrl_outclk_X13_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [2]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [2]),
	.Clk(\clk_25m~clkctrl_outclk_X12_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [3]),
	.Clk(\clk_25m~clkctrl_outclk_X3_Y7_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X3_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .coord_x = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [4]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [4]),
	.Clk(\clk_25m~clkctrl_outclk_X13_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [5]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [5]),
	.Clk(\clk_25m~clkctrl_outclk_X12_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [6]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [6]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [7]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [7]),
	.Clk(\clk_25m~clkctrl_outclk_X13_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [8]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [8]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [9]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [9]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [0]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [0]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [0]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(SyncReset_X16_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y12_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~5_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .mask = 16'h6FF6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [10]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y14_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [1]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [1]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [1]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(SyncReset_X16_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y12_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|data_wire[2]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .mask = 16'h0FF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [2]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [5]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [2]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y12_SIG ),
	.SyncReset(SyncReset_X16_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y12_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~3_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .mask = 16'h7DBE;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [3]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3]),
	.Clk(\clk_25m~clkctrl_outclk_X3_Y7_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X3_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .coord_x = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [7]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [4]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [4]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [7]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [4]),
	.Clk(\clk_25m~clkctrl_outclk_X13_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ),
	.SyncReset(SyncReset_X13_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y12_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~2_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .mask = 16'h7DBE;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [5]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [5]),
	.Clk(\clk_25m~clkctrl_outclk_X12_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ),
	.SyncReset(SyncReset_X12_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y13_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [6]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [6]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(SyncReset_X17_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X17_Y13_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~1_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .mask = 16'h6FF6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [7]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [7]),
	.Clk(\clk_25m~clkctrl_outclk_X13_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [8]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [8]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(SyncReset_X17_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X17_Y13_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .mask = 16'h6FF6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [9]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 (
	.A(\eth_udp_inst|ip_send_inst|read_data_req~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~5_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|data_wire[2]~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .mask = 16'hAAA8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|data_wire[2]~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~5_combout ),
	.C(\camera_if_inst|cam_hsync_r [1]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .mask = 16'hF0E0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~1_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~3_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~0_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .mask = 16'hFFFE;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .mask = 16'h0200;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .mask = 16'h0100;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .mask = 16'h0100;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .mask = 16'h0400;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .mask = 16'h0200;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .mask = 16'hC000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X13_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~6_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .mask = 16'hA5A5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [10]),
	.Clk(\cam_pclk~input_o_X13_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .mask = 16'hD2D2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1]),
	.Clk(\cam_pclk~input_o_X13_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1]~8_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .mask = 16'h78F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.Clk(\cam_pclk~input_o_X12_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2]~7_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .mask = 16'hD2F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]),
	.Clk(\cam_pclk~input_o_X12_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3]~9_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .mask = 16'h3CF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4]),
	.Clk(\cam_pclk~input_o_X12_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4]~5_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .mask = 16'hD2F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.Clk(\cam_pclk~input_o_X12_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5]~6_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .mask = 16'h3C3C;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]),
	.Clk(\cam_pclk~input_o_X13_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6]~3_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .mask = 16'h5AF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7]),
	.Clk(\cam_pclk~input_o_X13_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7]~4_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .mask = 16'hD2F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8]),
	.Clk(\cam_pclk~input_o_X13_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8]~1_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .mask = 16'h0FF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [9]),
	.Clk(\cam_pclk~input_o_X13_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9]~2_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .mask = 16'h7878;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X13_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~7_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .mask = 16'h6699;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0~q ),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X13_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~8_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .mask = 16'h9669;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1~q ),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X13_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~9_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [10]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [9]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2~q ),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X13_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~10_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .mask = 16'h9696;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .mask = 16'h3333;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(SyncReset_X16_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y13_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [12]),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [9]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [11]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(SyncReset_X16_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y13_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [11]),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [11]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .mask = 16'h5A5A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [10]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [12]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [12]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [1]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(SyncReset_X16_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y13_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y13_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(SyncReset_X14_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y13_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [0]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [0]),
	.Clk(\cam_pclk~input_o_X14_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [10]),
	.Clk(\cam_pclk~input_o_X16_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [1]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [1]),
	.Clk(\cam_pclk~input_o_X14_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(SyncReset_X14_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y13_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [2]),
	.Clk(\cam_pclk~input_o_X12_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ),
	.SyncReset(SyncReset_X12_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y13_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [3]),
	.Clk(\cam_pclk~input_o_X14_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [4]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [4]),
	.Clk(\cam_pclk~input_o_X13_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ),
	.SyncReset(SyncReset_X13_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y12_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [5]),
	.Clk(\cam_pclk~input_o_X12_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ),
	.SyncReset(SyncReset_X12_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y13_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [6]),
	.Clk(\cam_pclk~input_o_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [7]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [7]),
	.Clk(\cam_pclk~input_o_X13_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ),
	.SyncReset(SyncReset_X13_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y12_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [8]),
	.Clk(\cam_pclk~input_o_X16_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(SyncReset_X16_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y13_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [9]),
	.Clk(\cam_pclk~input_o_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [3]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [0]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [0]),
	.Clk(\cam_pclk~input_o_X14_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(SyncReset_X14_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y13_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~5_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .mask = 16'h7BDE;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [10]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [10]),
	.Clk(\cam_pclk~input_o_X16_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [1]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [1]),
	.Clk(\cam_pclk~input_o_X14_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(SyncReset_X14_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y13_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|data_wire[2]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .mask = 16'h3C3C;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [5]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [2]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [2]),
	.Clk(\cam_pclk~input_o_X12_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ),
	.SyncReset(SyncReset_X12_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y13_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~3_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .mask = 16'h6FF6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [3]),
	.Clk(\cam_pclk~input_o_X14_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [7]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [4]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [4]),
	.Clk(\cam_pclk~input_o_X13_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ),
	.SyncReset(SyncReset_X13_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y12_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~2_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .mask = 16'h6FF6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [5]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [5]),
	.Clk(\cam_pclk~input_o_X12_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [9]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [11]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [6]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [6]),
	.Clk(\cam_pclk~input_o_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(SyncReset_X17_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X17_Y13_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~1_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .mask = 16'h9FF9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [7]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [7]),
	.Clk(\cam_pclk~input_o_X13_Y12_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .coord_y = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [12]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [10]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [8]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [8]),
	.Clk(\cam_pclk~input_o_X16_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y13_SIG ),
	.SyncReset(SyncReset_X16_Y13_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y13_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .coord_y = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .mask = 16'h9FF9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [9]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [9]),
	.Clk(\cam_pclk~input_o_X17_Y13_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .coord_y = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .CarryEnb = 1'b1;

alta_dio \e_rx[0]~input (
	.padio(e_rx[0]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\e_rx[0]~input_o ),
	.regout());
defparam \e_rx[0]~input .coord_x = 49;
defparam \e_rx[0]~input .coord_y = 19;
defparam \e_rx[0]~input .coord_z = 0;
defparam \e_rx[0]~input .IN_ASYNC_MODE = 1'b0;
defparam \e_rx[0]~input .IN_SYNC_MODE = 1'b0;
defparam \e_rx[0]~input .IN_POWERUP = 1'b0;
defparam \e_rx[0]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \e_rx[0]~input .IN_SYNC_DISABLE = 1'b0;
defparam \e_rx[0]~input .OUT_REG_MODE = 1'b0;
defparam \e_rx[0]~input .OUT_ASYNC_MODE = 1'b0;
defparam \e_rx[0]~input .OUT_SYNC_MODE = 1'b0;
defparam \e_rx[0]~input .OUT_POWERUP = 1'b0;
defparam \e_rx[0]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_rx[0]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_rx[0]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \e_rx[0]~input .OUT_DDIO = 1'b0;
defparam \e_rx[0]~input .OE_REG_MODE = 1'b0;
defparam \e_rx[0]~input .OE_ASYNC_MODE = 1'b0;
defparam \e_rx[0]~input .OE_SYNC_MODE = 1'b0;
defparam \e_rx[0]~input .OE_POWERUP = 1'b0;
defparam \e_rx[0]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \e_rx[0]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \e_rx[0]~input .OE_SYNC_DISABLE = 1'b0;
defparam \e_rx[0]~input .OE_DDIO = 1'b0;
defparam \e_rx[0]~input .CFG_TRI_INPUT = 1'b0;
defparam \e_rx[0]~input .CFG_PULL_UP = 1'b0;
defparam \e_rx[0]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \e_rx[0]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_rx[0]~input .CFG_PDRV = 7'b0011010;
defparam \e_rx[0]~input .CFG_NDRV = 7'b0011000;
defparam \e_rx[0]~input .CFG_KEEP = 2'b00;
defparam \e_rx[0]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_rx[0]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_rx[0]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_rx[0]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \e_rx[0]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_rx[0]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_rx[0]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_rx[0]~input .CFG_OSCDIV = 2'b00;
defparam \e_rx[0]~input .CFG_ROCTUSR = 1'b0;
defparam \e_rx[0]~input .CFG_SEL_CUA = 1'b0;
defparam \e_rx[0]~input .CFG_ROCT_EN = 1'b0;
defparam \e_rx[0]~input .INPUT_ONLY = 1'b0;
defparam \e_rx[0]~input .DPCLK_DELAY = 4'b0000;
defparam \e_rx[0]~input .OUT_DELAY = 1'b0;
defparam \e_rx[0]~input .IN_DATA_DELAY = 3'b000;
defparam \e_rx[0]~input .IN_REG_DELAY = 3'b000;

alta_dio \e_rx[1]~input (
	.padio(e_rx[1]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\e_rx[1]~input_o ),
	.regout());
defparam \e_rx[1]~input .coord_x = 49;
defparam \e_rx[1]~input .coord_y = 20;
defparam \e_rx[1]~input .coord_z = 2;
defparam \e_rx[1]~input .IN_ASYNC_MODE = 1'b0;
defparam \e_rx[1]~input .IN_SYNC_MODE = 1'b0;
defparam \e_rx[1]~input .IN_POWERUP = 1'b0;
defparam \e_rx[1]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \e_rx[1]~input .IN_SYNC_DISABLE = 1'b0;
defparam \e_rx[1]~input .OUT_REG_MODE = 1'b0;
defparam \e_rx[1]~input .OUT_ASYNC_MODE = 1'b0;
defparam \e_rx[1]~input .OUT_SYNC_MODE = 1'b0;
defparam \e_rx[1]~input .OUT_POWERUP = 1'b0;
defparam \e_rx[1]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_rx[1]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_rx[1]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \e_rx[1]~input .OUT_DDIO = 1'b0;
defparam \e_rx[1]~input .OE_REG_MODE = 1'b0;
defparam \e_rx[1]~input .OE_ASYNC_MODE = 1'b0;
defparam \e_rx[1]~input .OE_SYNC_MODE = 1'b0;
defparam \e_rx[1]~input .OE_POWERUP = 1'b0;
defparam \e_rx[1]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \e_rx[1]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \e_rx[1]~input .OE_SYNC_DISABLE = 1'b0;
defparam \e_rx[1]~input .OE_DDIO = 1'b0;
defparam \e_rx[1]~input .CFG_TRI_INPUT = 1'b0;
defparam \e_rx[1]~input .CFG_PULL_UP = 1'b0;
defparam \e_rx[1]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \e_rx[1]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_rx[1]~input .CFG_PDRV = 7'b0011010;
defparam \e_rx[1]~input .CFG_NDRV = 7'b0011000;
defparam \e_rx[1]~input .CFG_KEEP = 2'b00;
defparam \e_rx[1]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_rx[1]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_rx[1]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_rx[1]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \e_rx[1]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_rx[1]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_rx[1]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_rx[1]~input .CFG_OSCDIV = 2'b00;
defparam \e_rx[1]~input .CFG_ROCTUSR = 1'b0;
defparam \e_rx[1]~input .CFG_SEL_CUA = 1'b0;
defparam \e_rx[1]~input .CFG_ROCT_EN = 1'b0;
defparam \e_rx[1]~input .INPUT_ONLY = 1'b0;
defparam \e_rx[1]~input .DPCLK_DELAY = 4'b0000;
defparam \e_rx[1]~input .OUT_DELAY = 1'b0;
defparam \e_rx[1]~input .IN_DATA_DELAY = 3'b000;
defparam \e_rx[1]~input .IN_REG_DELAY = 3'b000;

alta_dio \e_rxclk~input (
	.padio(e_rxclk),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\e_rxclk~input_o ),
	.regout());
defparam \e_rxclk~input .coord_x = 49;
defparam \e_rxclk~input .coord_y = 27;
defparam \e_rxclk~input .coord_z = 2;
defparam \e_rxclk~input .IN_ASYNC_MODE = 1'b0;
defparam \e_rxclk~input .IN_SYNC_MODE = 1'b0;
defparam \e_rxclk~input .IN_POWERUP = 1'b0;
defparam \e_rxclk~input .IN_ASYNC_DISABLE = 1'b0;
defparam \e_rxclk~input .IN_SYNC_DISABLE = 1'b0;
defparam \e_rxclk~input .OUT_REG_MODE = 1'b0;
defparam \e_rxclk~input .OUT_ASYNC_MODE = 1'b0;
defparam \e_rxclk~input .OUT_SYNC_MODE = 1'b0;
defparam \e_rxclk~input .OUT_POWERUP = 1'b0;
defparam \e_rxclk~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_rxclk~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_rxclk~input .OUT_SYNC_DISABLE = 1'b0;
defparam \e_rxclk~input .OUT_DDIO = 1'b0;
defparam \e_rxclk~input .OE_REG_MODE = 1'b0;
defparam \e_rxclk~input .OE_ASYNC_MODE = 1'b0;
defparam \e_rxclk~input .OE_SYNC_MODE = 1'b0;
defparam \e_rxclk~input .OE_POWERUP = 1'b0;
defparam \e_rxclk~input .OE_CLKEN_DISABLE = 1'b0;
defparam \e_rxclk~input .OE_ASYNC_DISABLE = 1'b0;
defparam \e_rxclk~input .OE_SYNC_DISABLE = 1'b0;
defparam \e_rxclk~input .OE_DDIO = 1'b0;
defparam \e_rxclk~input .CFG_TRI_INPUT = 1'b0;
defparam \e_rxclk~input .CFG_PULL_UP = 1'b0;
defparam \e_rxclk~input .CFG_OPEN_DRAIN = 1'b0;
defparam \e_rxclk~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_rxclk~input .CFG_PDRV = 7'b0011010;
defparam \e_rxclk~input .CFG_NDRV = 7'b0011000;
defparam \e_rxclk~input .CFG_KEEP = 2'b00;
defparam \e_rxclk~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_rxclk~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_rxclk~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_rxclk~input .CFG_LVDS_IN_EN = 1'b0;
defparam \e_rxclk~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_rxclk~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_rxclk~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_rxclk~input .CFG_OSCDIV = 2'b00;
defparam \e_rxclk~input .CFG_ROCTUSR = 1'b0;
defparam \e_rxclk~input .CFG_SEL_CUA = 1'b0;
defparam \e_rxclk~input .CFG_ROCT_EN = 1'b0;
defparam \e_rxclk~input .INPUT_ONLY = 1'b0;
defparam \e_rxclk~input .DPCLK_DELAY = 4'b0000;
defparam \e_rxclk~input .OUT_DELAY = 1'b0;
defparam \e_rxclk~input .IN_DATA_DELAY = 3'b000;
defparam \e_rxclk~input .IN_REG_DELAY = 3'b000;

alta_dio \e_rxdv~input (
	.padio(e_rxdv),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\e_rxdv~input_o ),
	.regout());
defparam \e_rxdv~input .coord_x = 49;
defparam \e_rxdv~input .coord_y = 19;
defparam \e_rxdv~input .coord_z = 3;
defparam \e_rxdv~input .IN_ASYNC_MODE = 1'b0;
defparam \e_rxdv~input .IN_SYNC_MODE = 1'b0;
defparam \e_rxdv~input .IN_POWERUP = 1'b0;
defparam \e_rxdv~input .IN_ASYNC_DISABLE = 1'b0;
defparam \e_rxdv~input .IN_SYNC_DISABLE = 1'b0;
defparam \e_rxdv~input .OUT_REG_MODE = 1'b0;
defparam \e_rxdv~input .OUT_ASYNC_MODE = 1'b0;
defparam \e_rxdv~input .OUT_SYNC_MODE = 1'b0;
defparam \e_rxdv~input .OUT_POWERUP = 1'b0;
defparam \e_rxdv~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_rxdv~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_rxdv~input .OUT_SYNC_DISABLE = 1'b0;
defparam \e_rxdv~input .OUT_DDIO = 1'b0;
defparam \e_rxdv~input .OE_REG_MODE = 1'b0;
defparam \e_rxdv~input .OE_ASYNC_MODE = 1'b0;
defparam \e_rxdv~input .OE_SYNC_MODE = 1'b0;
defparam \e_rxdv~input .OE_POWERUP = 1'b0;
defparam \e_rxdv~input .OE_CLKEN_DISABLE = 1'b0;
defparam \e_rxdv~input .OE_ASYNC_DISABLE = 1'b0;
defparam \e_rxdv~input .OE_SYNC_DISABLE = 1'b0;
defparam \e_rxdv~input .OE_DDIO = 1'b0;
defparam \e_rxdv~input .CFG_TRI_INPUT = 1'b0;
defparam \e_rxdv~input .CFG_PULL_UP = 1'b0;
defparam \e_rxdv~input .CFG_OPEN_DRAIN = 1'b0;
defparam \e_rxdv~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_rxdv~input .CFG_PDRV = 7'b0011010;
defparam \e_rxdv~input .CFG_NDRV = 7'b0011000;
defparam \e_rxdv~input .CFG_KEEP = 2'b00;
defparam \e_rxdv~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_rxdv~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_rxdv~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_rxdv~input .CFG_LVDS_IN_EN = 1'b0;
defparam \e_rxdv~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_rxdv~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_rxdv~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_rxdv~input .CFG_OSCDIV = 2'b00;
defparam \e_rxdv~input .CFG_ROCTUSR = 1'b0;
defparam \e_rxdv~input .CFG_SEL_CUA = 1'b0;
defparam \e_rxdv~input .CFG_ROCT_EN = 1'b0;
defparam \e_rxdv~input .INPUT_ONLY = 1'b0;
defparam \e_rxdv~input .DPCLK_DELAY = 4'b0000;
defparam \e_rxdv~input .OUT_DELAY = 1'b0;
defparam \e_rxdv~input .IN_DATA_DELAY = 3'b000;
defparam \e_rxdv~input .IN_REG_DELAY = 3'b000;

alta_dio \e_rxer~input (
	.padio(e_rxer),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\e_rxer~input_o ),
	.regout());
defparam \e_rxer~input .coord_x = 49;
defparam \e_rxer~input .coord_y = 19;
defparam \e_rxer~input .coord_z = 1;
defparam \e_rxer~input .IN_ASYNC_MODE = 1'b0;
defparam \e_rxer~input .IN_SYNC_MODE = 1'b0;
defparam \e_rxer~input .IN_POWERUP = 1'b0;
defparam \e_rxer~input .IN_ASYNC_DISABLE = 1'b0;
defparam \e_rxer~input .IN_SYNC_DISABLE = 1'b0;
defparam \e_rxer~input .OUT_REG_MODE = 1'b0;
defparam \e_rxer~input .OUT_ASYNC_MODE = 1'b0;
defparam \e_rxer~input .OUT_SYNC_MODE = 1'b0;
defparam \e_rxer~input .OUT_POWERUP = 1'b0;
defparam \e_rxer~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_rxer~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_rxer~input .OUT_SYNC_DISABLE = 1'b0;
defparam \e_rxer~input .OUT_DDIO = 1'b0;
defparam \e_rxer~input .OE_REG_MODE = 1'b0;
defparam \e_rxer~input .OE_ASYNC_MODE = 1'b0;
defparam \e_rxer~input .OE_SYNC_MODE = 1'b0;
defparam \e_rxer~input .OE_POWERUP = 1'b0;
defparam \e_rxer~input .OE_CLKEN_DISABLE = 1'b0;
defparam \e_rxer~input .OE_ASYNC_DISABLE = 1'b0;
defparam \e_rxer~input .OE_SYNC_DISABLE = 1'b0;
defparam \e_rxer~input .OE_DDIO = 1'b0;
defparam \e_rxer~input .CFG_TRI_INPUT = 1'b0;
defparam \e_rxer~input .CFG_PULL_UP = 1'b0;
defparam \e_rxer~input .CFG_OPEN_DRAIN = 1'b0;
defparam \e_rxer~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_rxer~input .CFG_PDRV = 7'b0011010;
defparam \e_rxer~input .CFG_NDRV = 7'b0011000;
defparam \e_rxer~input .CFG_KEEP = 2'b00;
defparam \e_rxer~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_rxer~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_rxer~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_rxer~input .CFG_LVDS_IN_EN = 1'b0;
defparam \e_rxer~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_rxer~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_rxer~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_rxer~input .CFG_OSCDIV = 2'b00;
defparam \e_rxer~input .CFG_ROCTUSR = 1'b0;
defparam \e_rxer~input .CFG_SEL_CUA = 1'b0;
defparam \e_rxer~input .CFG_ROCT_EN = 1'b0;
defparam \e_rxer~input .INPUT_ONLY = 1'b0;
defparam \e_rxer~input .DPCLK_DELAY = 4'b0000;
defparam \e_rxer~input .OUT_DELAY = 1'b0;
defparam \e_rxer~input .IN_DATA_DELAY = 3'b000;
defparam \e_rxer~input .IN_REG_DELAY = 3'b000;

alta_dio \e_tx[0]~output (
	.padio(e_tx[0]),
	.datain(\mii_to_rmii_inst|eth_tx_data [0]),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \e_tx[0]~output .coord_x = 49;
defparam \e_tx[0]~output .coord_y = 27;
defparam \e_tx[0]~output .coord_z = 1;
defparam \e_tx[0]~output .IN_ASYNC_MODE = 1'b0;
defparam \e_tx[0]~output .IN_SYNC_MODE = 1'b0;
defparam \e_tx[0]~output .IN_POWERUP = 1'b0;
defparam \e_tx[0]~output .IN_ASYNC_DISABLE = 1'b0;
defparam \e_tx[0]~output .IN_SYNC_DISABLE = 1'b0;
defparam \e_tx[0]~output .OUT_REG_MODE = 1'b0;
defparam \e_tx[0]~output .OUT_ASYNC_MODE = 1'b0;
defparam \e_tx[0]~output .OUT_SYNC_MODE = 1'b0;
defparam \e_tx[0]~output .OUT_POWERUP = 1'b0;
defparam \e_tx[0]~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_tx[0]~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_tx[0]~output .OUT_SYNC_DISABLE = 1'b0;
defparam \e_tx[0]~output .OUT_DDIO = 1'b0;
defparam \e_tx[0]~output .OE_REG_MODE = 1'b0;
defparam \e_tx[0]~output .OE_ASYNC_MODE = 1'b0;
defparam \e_tx[0]~output .OE_SYNC_MODE = 1'b0;
defparam \e_tx[0]~output .OE_POWERUP = 1'b0;
defparam \e_tx[0]~output .OE_CLKEN_DISABLE = 1'b0;
defparam \e_tx[0]~output .OE_ASYNC_DISABLE = 1'b0;
defparam \e_tx[0]~output .OE_SYNC_DISABLE = 1'b0;
defparam \e_tx[0]~output .OE_DDIO = 1'b0;
defparam \e_tx[0]~output .CFG_TRI_INPUT = 1'b0;
defparam \e_tx[0]~output .CFG_PULL_UP = 1'b0;
defparam \e_tx[0]~output .CFG_OPEN_DRAIN = 1'b0;
defparam \e_tx[0]~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_tx[0]~output .CFG_PDRV = 7'b0011010;
defparam \e_tx[0]~output .CFG_NDRV = 7'b0011000;
defparam \e_tx[0]~output .CFG_KEEP = 2'b00;
defparam \e_tx[0]~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_tx[0]~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_tx[0]~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_tx[0]~output .CFG_LVDS_IN_EN = 1'b0;
defparam \e_tx[0]~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_tx[0]~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_tx[0]~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_tx[0]~output .CFG_OSCDIV = 2'b00;
defparam \e_tx[0]~output .CFG_ROCTUSR = 1'b0;
defparam \e_tx[0]~output .CFG_SEL_CUA = 1'b0;
defparam \e_tx[0]~output .CFG_ROCT_EN = 1'b0;
defparam \e_tx[0]~output .INPUT_ONLY = 1'b0;
defparam \e_tx[0]~output .DPCLK_DELAY = 4'b0000;
defparam \e_tx[0]~output .OUT_DELAY = 1'b0;
defparam \e_tx[0]~output .IN_DATA_DELAY = 3'b000;
defparam \e_tx[0]~output .IN_REG_DELAY = 3'b000;

alta_dio \e_tx[1]~output (
	.padio(e_tx[1]),
	.datain(\mii_to_rmii_inst|eth_tx_data [1]),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \e_tx[1]~output .coord_x = 44;
defparam \e_tx[1]~output .coord_y = 29;
defparam \e_tx[1]~output .coord_z = 2;
defparam \e_tx[1]~output .IN_ASYNC_MODE = 1'b0;
defparam \e_tx[1]~output .IN_SYNC_MODE = 1'b0;
defparam \e_tx[1]~output .IN_POWERUP = 1'b0;
defparam \e_tx[1]~output .IN_ASYNC_DISABLE = 1'b0;
defparam \e_tx[1]~output .IN_SYNC_DISABLE = 1'b0;
defparam \e_tx[1]~output .OUT_REG_MODE = 1'b0;
defparam \e_tx[1]~output .OUT_ASYNC_MODE = 1'b0;
defparam \e_tx[1]~output .OUT_SYNC_MODE = 1'b0;
defparam \e_tx[1]~output .OUT_POWERUP = 1'b0;
defparam \e_tx[1]~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_tx[1]~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_tx[1]~output .OUT_SYNC_DISABLE = 1'b0;
defparam \e_tx[1]~output .OUT_DDIO = 1'b0;
defparam \e_tx[1]~output .OE_REG_MODE = 1'b0;
defparam \e_tx[1]~output .OE_ASYNC_MODE = 1'b0;
defparam \e_tx[1]~output .OE_SYNC_MODE = 1'b0;
defparam \e_tx[1]~output .OE_POWERUP = 1'b0;
defparam \e_tx[1]~output .OE_CLKEN_DISABLE = 1'b0;
defparam \e_tx[1]~output .OE_ASYNC_DISABLE = 1'b0;
defparam \e_tx[1]~output .OE_SYNC_DISABLE = 1'b0;
defparam \e_tx[1]~output .OE_DDIO = 1'b0;
defparam \e_tx[1]~output .CFG_TRI_INPUT = 1'b0;
defparam \e_tx[1]~output .CFG_PULL_UP = 1'b0;
defparam \e_tx[1]~output .CFG_OPEN_DRAIN = 1'b0;
defparam \e_tx[1]~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_tx[1]~output .CFG_PDRV = 7'b0011010;
defparam \e_tx[1]~output .CFG_NDRV = 7'b0011000;
defparam \e_tx[1]~output .CFG_KEEP = 2'b00;
defparam \e_tx[1]~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_tx[1]~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_tx[1]~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_tx[1]~output .CFG_LVDS_IN_EN = 1'b0;
defparam \e_tx[1]~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_tx[1]~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_tx[1]~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_tx[1]~output .CFG_OSCDIV = 2'b00;
defparam \e_tx[1]~output .CFG_ROCTUSR = 1'b0;
defparam \e_tx[1]~output .CFG_SEL_CUA = 1'b0;
defparam \e_tx[1]~output .CFG_ROCT_EN = 1'b0;
defparam \e_tx[1]~output .INPUT_ONLY = 1'b0;
defparam \e_tx[1]~output .DPCLK_DELAY = 4'b0000;
defparam \e_tx[1]~output .OUT_DELAY = 1'b0;
defparam \e_tx[1]~output .IN_DATA_DELAY = 3'b000;
defparam \e_tx[1]~output .IN_REG_DELAY = 3'b000;

alta_dio \e_txen~output (
	.padio(e_txen),
	.datain(\mii_to_rmii_inst|eth_tx_dv~q ),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \e_txen~output .coord_x = 43;
defparam \e_txen~output .coord_y = 29;
defparam \e_txen~output .coord_z = 1;
defparam \e_txen~output .IN_ASYNC_MODE = 1'b0;
defparam \e_txen~output .IN_SYNC_MODE = 1'b0;
defparam \e_txen~output .IN_POWERUP = 1'b0;
defparam \e_txen~output .IN_ASYNC_DISABLE = 1'b0;
defparam \e_txen~output .IN_SYNC_DISABLE = 1'b0;
defparam \e_txen~output .OUT_REG_MODE = 1'b0;
defparam \e_txen~output .OUT_ASYNC_MODE = 1'b0;
defparam \e_txen~output .OUT_SYNC_MODE = 1'b0;
defparam \e_txen~output .OUT_POWERUP = 1'b0;
defparam \e_txen~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_txen~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_txen~output .OUT_SYNC_DISABLE = 1'b0;
defparam \e_txen~output .OUT_DDIO = 1'b0;
defparam \e_txen~output .OE_REG_MODE = 1'b0;
defparam \e_txen~output .OE_ASYNC_MODE = 1'b0;
defparam \e_txen~output .OE_SYNC_MODE = 1'b0;
defparam \e_txen~output .OE_POWERUP = 1'b0;
defparam \e_txen~output .OE_CLKEN_DISABLE = 1'b0;
defparam \e_txen~output .OE_ASYNC_DISABLE = 1'b0;
defparam \e_txen~output .OE_SYNC_DISABLE = 1'b0;
defparam \e_txen~output .OE_DDIO = 1'b0;
defparam \e_txen~output .CFG_TRI_INPUT = 1'b0;
defparam \e_txen~output .CFG_PULL_UP = 1'b0;
defparam \e_txen~output .CFG_OPEN_DRAIN = 1'b0;
defparam \e_txen~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_txen~output .CFG_PDRV = 7'b0011010;
defparam \e_txen~output .CFG_NDRV = 7'b0011000;
defparam \e_txen~output .CFG_KEEP = 2'b00;
defparam \e_txen~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_txen~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_txen~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_txen~output .CFG_LVDS_IN_EN = 1'b0;
defparam \e_txen~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_txen~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_txen~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_txen~output .CFG_OSCDIV = 2'b00;
defparam \e_txen~output .CFG_ROCTUSR = 1'b0;
defparam \e_txen~output .CFG_SEL_CUA = 1'b0;
defparam \e_txen~output .CFG_ROCT_EN = 1'b0;
defparam \e_txen~output .INPUT_ONLY = 1'b0;
defparam \e_txen~output .DPCLK_DELAY = 4'b0000;
defparam \e_txen~output .OUT_DELAY = 1'b0;
defparam \e_txen~output .IN_DATA_DELAY = 3'b000;
defparam \e_txen~output .IN_REG_DELAY = 3'b000;

alta_slice \eth_udp_inst|crc32_inst|crc_data[0] (
	.A(vcc),
	.B(\eth_udp_inst|crc32_inst|crc_data [28]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [0]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~25_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [0]));
defparam \eth_udp_inst|crc32_inst|crc_data[0] .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .coord_z = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .mask = 16'h003C;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[10] (
	.A(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.B(\eth_udp_inst|crc32_inst|crc_data [6]),
	.C(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [10]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~30_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [10]));
defparam \eth_udp_inst|crc32_inst|crc_data[10] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .coord_z = 7;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[11] (
	.A(\eth_udp_inst|crc32_inst|crc_next~5_combout ),
	.B(\eth_udp_inst|crc32_inst|crc_data [7]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [11]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~16_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [11]));
defparam \eth_udp_inst|crc32_inst|crc_data[11] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .coord_z = 15;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .mask = 16'h0066;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[12] (
	.A(\eth_udp_inst|crc32_inst|crc_next~2_combout ),
	.B(\eth_udp_inst|crc32_inst|crc_data [8]),
	.C(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [12]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~24_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [12]));
defparam \eth_udp_inst|crc32_inst|crc_data[12] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .coord_z = 1;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[13] (
	.A(\eth_udp_inst|crc32_inst|crc_data [9]),
	.B(\eth_udp_inst|crc32_inst|crc_next~6_combout ),
	.C(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [13]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~11_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [13]));
defparam \eth_udp_inst|crc32_inst|crc_data[13] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .coord_z = 11;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[14] (
	.A(vcc),
	.B(\eth_udp_inst|crc32_inst|crc_data [10]),
	.C(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [14]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~32_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [14]));
defparam \eth_udp_inst|crc32_inst|crc_data[14] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .coord_z = 15;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .mask = 16'h003C;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[15] (
	.A(\eth_udp_inst|crc32_inst|crc_data [11]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.C(\eth_udp_inst|crc32_inst|crc_data [31]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [15]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~18_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [15]));
defparam \eth_udp_inst|crc32_inst|crc_data[15] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .coord_z = 8;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[16] (
	.A(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.B(\eth_udp_inst|crc32_inst|crc_data [28]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.D(\eth_udp_inst|crc32_inst|crc_data [12]),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [16]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~29_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [16]));
defparam \eth_udp_inst|crc32_inst|crc_data[16] .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .coord_z = 7;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .mask = 16'h1441;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[17] (
	.A(\eth_udp_inst|crc32_inst|crc_data [29]),
	.B(\eth_udp_inst|crc32_inst|crc_data [13]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [17]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~15_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [17]));
defparam \eth_udp_inst|crc32_inst|crc_data[17] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .coord_z = 10;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[18] (
	.A(\eth_udp_inst|crc32_inst|crc_data [14]),
	.B(\eth_udp_inst|crc32_inst|crc_data [30]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [18]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~35_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [18]));
defparam \eth_udp_inst|crc32_inst|crc_data[18] .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .coord_z = 3;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[19] (
	.A(\eth_udp_inst|crc32_inst|crc_data [31]),
	.B(\eth_udp_inst|crc32_inst|crc_data [15]),
	.C(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [19]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~21_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [19]));
defparam \eth_udp_inst|crc32_inst|crc_data[19] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .coord_z = 2;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .mask = 16'h0609;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[1] (
	.A(\eth_udp_inst|crc32_inst|crc_data [29]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.C(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [1]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~38_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [1]));
defparam \eth_udp_inst|crc32_inst|crc_data[1] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .coord_z = 12;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[20] (
	.A(vcc),
	.B(\eth_udp_inst|crc32_inst|crc_data [16]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [20]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~26_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [20]));
defparam \eth_udp_inst|crc32_inst|crc_data[20] .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .coord_z = 10;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .mask = 16'h00CC;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[21] (
	.A(vcc),
	.B(\eth_udp_inst|crc32_inst|crc_data [17]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [21]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~12_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [21]));
defparam \eth_udp_inst|crc32_inst|crc_data[21] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .coord_z = 0;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .mask = 16'h00CC;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[22] (
	.A(\eth_udp_inst|crc32_inst|crc_data [18]),
	.B(\eth_udp_inst|crc32_inst|crc_data [28]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [22]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~33_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [22]));
defparam \eth_udp_inst|crc32_inst|crc_data[22] .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .coord_z = 15;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[23] (
	.A(\eth_udp_inst|crc32_inst|crc_data [19]),
	.B(\eth_udp_inst|crc32_inst|crc_next~6_combout ),
	.C(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [23]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~19_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [23]));
defparam \eth_udp_inst|crc32_inst|crc_data[23] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .coord_z = 13;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .mask = 16'h0096;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[24] (
	.A(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.B(\eth_udp_inst|crc32_inst|crc_data [20]),
	.C(vcc),
	.D(\eth_udp_inst|crc32_inst|crc_next~2_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [24]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~27_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [24]));
defparam \eth_udp_inst|crc32_inst|crc_data[24] .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .coord_z = 5;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .mask = 16'h1144;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[25] (
	.A(\eth_udp_inst|crc32_inst|crc_data [21]),
	.B(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [25]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~13_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [25]));
defparam \eth_udp_inst|crc32_inst|crc_data[25] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .coord_z = 6;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .mask = 16'h0066;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[26] (
	.A(\eth_udp_inst|crc32_inst|crc_data [22]),
	.B(\eth_udp_inst|crc32_inst|crc_next~3_combout ),
	.C(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [26]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~34_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [26]));
defparam \eth_udp_inst|crc32_inst|crc_data[26] .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .coord_z = 1;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .mask = 16'h0096;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[27] (
	.A(\eth_udp_inst|crc32_inst|crc_data [29]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.C(\eth_udp_inst|crc32_inst|crc_data [23]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [27]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~20_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [27]));
defparam \eth_udp_inst|crc32_inst|crc_data[27] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .coord_z = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[28] (
	.A(\eth_udp_inst|crc32_inst|crc_data [24]),
	.B(\eth_udp_inst|crc32_inst|crc_data [30]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [28]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~37_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [28]));
defparam \eth_udp_inst|crc32_inst|crc_data[28] .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .coord_z = 14;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[29] (
	.A(\eth_udp_inst|crc32_inst|crc_data [25]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.C(\eth_udp_inst|crc32_inst|crc_data [31]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [29]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~36_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [29]));
defparam \eth_udp_inst|crc32_inst|crc_data[29] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .coord_z = 11;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[2] (
	.A(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.B(\eth_udp_inst|crc32_inst|crc_data [28]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.D(\eth_udp_inst|crc32_inst|crc_next~2_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [2]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~40_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [2]));
defparam \eth_udp_inst|crc32_inst|crc_data[2] .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .coord_z = 6;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .mask = 16'h4114;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[30] (
	.A(\eth_udp_inst|crc32_inst|crc_data [26]),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [30]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~28_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [30]));
defparam \eth_udp_inst|crc32_inst|crc_data[30] .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .coord_z = 8;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .mask = 16'h00AA;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[31] (
	.A(vcc),
	.B(\eth_udp_inst|crc32_inst|crc_data [27]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [31]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~14_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [31]));
defparam \eth_udp_inst|crc32_inst|crc_data[31] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .coord_z = 3;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .mask = 16'h00CC;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[3] (
	.A(\eth_udp_inst|crc32_inst|crc_data [29]),
	.B(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [3]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~39_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [3]));
defparam \eth_udp_inst|crc32_inst|crc_data[3] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .coord_z = 1;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .mask = 16'h0096;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[4] (
	.A(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.B(\eth_udp_inst|crc32_inst|crc_data [0]),
	.C(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [4]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~23_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [4]));
defparam \eth_udp_inst|crc32_inst|crc_data[4] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .coord_z = 12;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[5] (
	.A(\eth_udp_inst|crc32_inst|crc_next~5_combout ),
	.B(vcc),
	.C(\eth_udp_inst|crc32_inst|crc_data [1]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [5]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~10_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [5]));
defparam \eth_udp_inst|crc32_inst|crc_data[5] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .coord_z = 6;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .mask = 16'h005A;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[6] (
	.A(\eth_udp_inst|crc32_inst|crc_data [2]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.D(\eth_udp_inst|crc32_inst|crc_next~2_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [6]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~31_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [6]));
defparam \eth_udp_inst|crc32_inst|crc_data[6] .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .coord_z = 4;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .mask = 16'h050A;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[7] (
	.A(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.B(\eth_udp_inst|crc32_inst|crc_data [3]),
	.C(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.D(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [7]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~17_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [7]));
defparam \eth_udp_inst|crc32_inst|crc_data[7] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .coord_z = 7;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .mask = 16'h0609;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[8] (
	.A(\eth_udp_inst|crc32_inst|crc_next~5_combout ),
	.B(\eth_udp_inst|crc32_inst|crc_data [4]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [8]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~22_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [8]));
defparam \eth_udp_inst|crc32_inst|crc_data[8] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .coord_z = 2;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .mask = 16'h0066;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[9] (
	.A(\eth_udp_inst|crc32_inst|crc_data [5]),
	.B(vcc),
	.C(\eth_udp_inst|crc32_inst|crc_next~2_combout ),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [9]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[28]~9_combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~8_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [9]));
defparam \eth_udp_inst|crc32_inst|crc_data[9] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .coord_z = 3;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .mask = 16'h005A;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next[28]~1 (
	.A(\eth_udp_inst|crc32_inst|crc_data [24]),
	.B(\eth_udp_inst|crc32_inst|crc_data [30]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.D(\eth_udp_inst|ip_send_inst|crc_en~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next[28]~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .coord_z = 2;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .mask = 16'h9600;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next[29]~0 (
	.A(\eth_udp_inst|crc32_inst|crc_data [31]),
	.B(\eth_udp_inst|crc32_inst|crc_data [25]),
	.C(\eth_udp_inst|ip_send_inst|crc_en~q ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next[29]~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .coord_z = 12;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .mask = 16'h9060;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next~2 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.B(\eth_udp_inst|crc32_inst|crc_data [30]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.D(\eth_udp_inst|crc32_inst|crc_data [29]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next~2 .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .coord_z = 9;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .mask = 16'h6996;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next~3 (
	.A(\eth_udp_inst|crc32_inst|crc_data [31]),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next~3 .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .coord_z = 8;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .mask = 16'h55AA;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next~4 (
	.A(vcc),
	.B(\eth_udp_inst|crc32_inst|crc_data [28]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next~4 .coord_x = 19;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .coord_z = 12;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .mask = 16'h3C3C;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next~5 (
	.A(\eth_udp_inst|crc32_inst|crc_data [29]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.C(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.D(\eth_udp_inst|crc32_inst|crc_next~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next~5_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next~5 .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .coord_y = 16;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .coord_z = 13;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .mask = 16'h9669;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next~6 (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.D(\eth_udp_inst|crc32_inst|crc_data [29]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next~6_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next~6 .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .coord_z = 6;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .mask = 16'h0FF0;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next~7 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.B(\eth_udp_inst|crc32_inst|crc_data [30]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.D(\eth_udp_inst|crc32_inst|crc_data [31]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next~7 .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .coord_y = 17;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .coord_z = 10;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .mask = 16'h6996;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add13~0 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|cnt_add [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .mask = 16'h6688;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~10 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~10 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~12 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~12 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~14 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~14 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~16 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [8]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~16 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~18 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [9]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~18 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~2 (
	.A(\eth_udp_inst|ip_send_inst|cnt_add [1]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~2 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~20 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [10]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~20 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~22 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [11]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~22 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~24 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [12]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~24 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~26 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [13]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~26 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~28 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [14]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~29 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~28 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~30 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [15]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~29 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~30_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~30 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .mask = 16'h3C3C;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add13~4 (
	.A(\eth_udp_inst|ip_send_inst|cnt_add [2]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~4 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~6 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [3]),
	.B(\eth_udp_inst|ip_send_inst|cnt_add [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~6 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~8 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [4]),
	.B(\eth_udp_inst|ip_send_inst|cnt_add [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~8 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .mask = 16'h6688;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~10 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~10 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~12 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~12 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .mask = 16'h962B;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~14 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~14 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~16 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~16 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .mask = 16'h962B;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~18 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~18 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~2 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~2 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~20 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~20 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~22 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~22 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~24 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~24 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .mask = 16'h3CCF;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~26 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~26 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~28 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~28_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~28 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .mask = 16'h0F0F;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add2~4 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~4 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~6 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~6 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~8 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~8 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add3~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add2~24_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add3~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add3~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add3~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .mask = 16'h33CC;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add3~2 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add2~26_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add3~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add3~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add3~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add3~2 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add3~4 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|Add2~28_combout ),
	.Cin(\eth_udp_inst|ip_send_inst|Add3~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add3~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add3~4 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .mask = 16'hF00F;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add4~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .mask = 16'h6688;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~10 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][5]~q ),
	.B(\eth_udp_inst|ip_send_inst|Add2~6_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~10 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~12 (
	.A(\eth_udp_inst|ip_send_inst|Add2~8_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][6]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~12 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~14 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][7]~q ),
	.B(\eth_udp_inst|ip_send_inst|Add2~10_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~14 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~16 (
	.A(\eth_udp_inst|ip_send_inst|Add2~12_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~16 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~18 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][9]~q ),
	.B(\eth_udp_inst|ip_send_inst|Add2~14_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~18 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~2 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][1]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~2 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~20 (
	.A(\eth_udp_inst|ip_send_inst|Add2~16_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][10]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~20 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~22 (
	.A(\eth_udp_inst|ip_send_inst|Add2~18_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][11]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~22 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~24 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][12]~q ),
	.B(\eth_udp_inst|ip_send_inst|Add2~20_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~24 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~26 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][13]~q ),
	.B(\eth_udp_inst|ip_send_inst|Add2~22_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~26 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~28 (
	.A(\eth_udp_inst|ip_send_inst|Add3~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][14]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~29 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~28 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~30 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][15]~q ),
	.B(\eth_udp_inst|ip_send_inst|Add3~2_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~29 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~30_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~31 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~30 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~32 (
	.A(\eth_udp_inst|ip_send_inst|Add3~4_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~31 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~32_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~33 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~32 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~34 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~33 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~34_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~34 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .mask = 16'hF0F0;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add4~4 (
	.A(\eth_udp_inst|ip_send_inst|Add2~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][2]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~4 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~6 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][3]~q ),
	.B(\eth_udp_inst|ip_send_inst|Add2~2_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~6 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~8 (
	.A(\eth_udp_inst|ip_send_inst|Add2~4_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][4]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~8 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~0_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .mask = 16'h33CC;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~10 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~10_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~10 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~12 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~12_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~12 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~14 (
	.A(\eth_udp_inst|ip_send_inst|Add4~14_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~14 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~16 (
	.A(\eth_udp_inst|ip_send_inst|Add4~16_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~16 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~18 (
	.A(\eth_udp_inst|ip_send_inst|Add4~18_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~18 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~2 (
	.A(\eth_udp_inst|ip_send_inst|Add4~2_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~2 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~20 (
	.A(\eth_udp_inst|ip_send_inst|Add4~20_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~20 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~22 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~22_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~22 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~24 (
	.A(\eth_udp_inst|ip_send_inst|Add4~24_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~24 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~26 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~26_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~26 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~28 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~28_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~29 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~28 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .mask = 16'h3CCF;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~30 (
	.A(\eth_udp_inst|ip_send_inst|Add4~30_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~29 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~30_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~31 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~30 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~32 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~32_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~31 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~32_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~33 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~32 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~34 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~34_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~33 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~34_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~34 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .mask = 16'h3C3C;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add5~4 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~4_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~4 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~6 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~6_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~6 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~8 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~8_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~8 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .mask = 16'h3CCF;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~6_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~0 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .mask = 16'h33CC;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~10 (
	.A(\eth_udp_inst|ip_send_inst|Add5~16_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~10 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~12 (
	.A(\eth_udp_inst|ip_send_inst|Add5~18_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~12 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~14 (
	.A(\eth_udp_inst|ip_send_inst|Add5~20_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~14 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~16 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~22_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~16 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~18 (
	.A(\eth_udp_inst|ip_send_inst|Add5~24_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~18 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~2 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~8_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~2 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~20 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~26_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~20 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~22 (
	.A(\eth_udp_inst|ip_send_inst|Add5~28_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~22 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .mask = 16'hA505;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~24 (
	.A(\eth_udp_inst|ip_send_inst|Add5~30_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~24 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .mask = 16'h5AAF;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~26 (
	.A(\eth_udp_inst|ip_send_inst|Add5~32_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~26 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~28 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~34_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~28_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~28 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .mask = 16'hC3C3;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add6~4 (
	.A(\eth_udp_inst|ip_send_inst|Add5~10_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~4 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .mask = 16'h5AAF;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~6 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~12_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~6 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~8 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~14_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~8 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .mask = 16'h3CCF;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~2_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~0 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .mask = 16'h33CC;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~10 (
	.A(\eth_udp_inst|ip_send_inst|Add6~6_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~10 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~12 (
	.A(\eth_udp_inst|ip_send_inst|Add6~8_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~12 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~14 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~10_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~14 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .mask = 16'hC303;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~16 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~12_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~16 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .mask = 16'h3CCF;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~18 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~14_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~18 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~2 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~4_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~2 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~20 (
	.A(\eth_udp_inst|ip_send_inst|Add6~16_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~20 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~22 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~18_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~22 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~24 (
	.A(\eth_udp_inst|ip_send_inst|Add6~20_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~24 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~26 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~22_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~26 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~28 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~24_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~29 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~28 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~30 (
	.A(\eth_udp_inst|ip_send_inst|Add6~26_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~29 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~30_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~31 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~30 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~32 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|Add6~28_combout ),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~31 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~32_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~32 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .mask = 16'hF00F;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add7~4 (
	.A(\eth_udp_inst|ip_send_inst|Add6~0_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~4 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~6 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~2_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~6 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~8 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~4_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~8 .coord_x = 25;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~4_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~0 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .mask = 16'h33CC;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~10 (
	.A(\eth_udp_inst|ip_send_inst|Add7~14_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~10 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~12 (
	.A(\eth_udp_inst|ip_send_inst|Add7~16_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~12 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~14 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~18_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~14 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~16 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~20_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~16 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~18 (
	.A(\eth_udp_inst|ip_send_inst|Add7~22_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~18 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~2 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~6_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~2 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~20 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~24_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~20 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~22 (
	.A(\eth_udp_inst|ip_send_inst|Add7~26_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~22 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .mask = 16'hA505;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~24 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~28_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~24 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .mask = 16'h3CCF;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~26 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~30_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~26 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~28 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~32_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~29 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~28 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~30 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~29 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~30_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~30 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .mask = 16'hF0F0;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add8~4 (
	.A(\eth_udp_inst|ip_send_inst|Add7~8_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~4 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .mask = 16'h5AAF;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~6 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~10_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~6 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~8 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~12_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~8 .coord_x = 24;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .mask = 16'h3CCF;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~0_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .mask = 16'h33CC;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~10 (
	.A(\eth_udp_inst|ip_send_inst|Add8~4_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~10 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~12 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~6_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~12 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~14 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~8_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~14 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~16 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~10_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~16 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .mask = 16'h3CCF;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~18 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~12_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~18 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .mask = 16'hC303;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~2 (
	.A(\eth_udp_inst|ip_send_inst|Add7~0_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~2 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .mask = 16'hA505;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~20 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~14_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~20 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~22 (
	.A(\eth_udp_inst|ip_send_inst|Add8~16_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~22 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~24 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~18_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~24 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~26 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~20_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~26 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~28 (
	.A(\eth_udp_inst|ip_send_inst|Add8~22_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~29 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~28 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~30 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~24_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~29 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~30_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~31 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~30 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~32 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~26_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~31 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~32_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~33 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~32 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~34 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~28_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~33 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~34_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~35 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~34 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~36 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|Add8~30_combout ),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~35 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~36_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~36 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .mask = 16'hF00F;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add9~4 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~2_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~4 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~6 (
	.A(\eth_udp_inst|ip_send_inst|Add8~0_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~6 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~8 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~2_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~8 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Equal1~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .mask = 16'h0505;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal1~1 (
	.A(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|cnt [4]),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal1~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .mask = 16'h0002;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~0 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [9]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [10]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .mask = 16'h4488;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~1 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [3]),
	.C(\eth_udp_inst|ip_send_inst|data_cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|data_cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .coord_y = 20;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .mask = 16'h8000;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~2 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [4]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [5]),
	.C(\eth_udp_inst|ip_send_inst|data_cnt [6]),
	.D(\eth_udp_inst|ip_send_inst|data_cnt [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .coord_y = 19;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .mask = 16'h8000;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~3 (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Equal8~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|Equal8~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .mask = 16'hF000;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~4 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [13]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [11]),
	.C(\eth_udp_inst|ip_send_inst|data_cnt [12]),
	.D(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .mask = 16'h0180;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~5 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [8]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [15]),
	.C(\eth_udp_inst|ip_send_inst|data_cnt [14]),
	.D(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~5_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .mask = 16'h0180;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~6 (
	.A(\eth_udp_inst|ip_send_inst|Equal8~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|Equal8~4_combout ),
	.C(\eth_udp_inst|ip_send_inst|Equal8~5_combout ),
	.D(\eth_udp_inst|ip_send_inst|Equal8~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~6_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .mask = 16'h8000;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal9~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .mask = 16'h0011;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~0 (
	.A(\eth_udp_inst|ip_send_inst|Add13~26_combout ),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add13~30_combout ),
	.D(\eth_udp_inst|ip_send_inst|Add13~28_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .coord_y = 19;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .mask = 16'hFFFA;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~1 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add13~22_combout ),
	.C(\eth_udp_inst|ip_send_inst|Add13~24_combout ),
	.D(\eth_udp_inst|ip_send_inst|LessThan1~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .coord_y = 19;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .mask = 16'hFFFC;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~2 (
	.A(\eth_udp_inst|ip_send_inst|Add13~14_combout ),
	.B(\eth_udp_inst|ip_send_inst|Add13~12_combout ),
	.C(\eth_udp_inst|ip_send_inst|Add13~20_combout ),
	.D(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .mask = 16'h88FE;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~3 (
	.A(\eth_udp_inst|ip_send_inst|Add13~4_combout ),
	.B(\eth_udp_inst|ip_send_inst|data_len [10]),
	.C(\eth_udp_inst|ip_send_inst|Add13~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|Add13~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .mask = 16'hB332;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~4 (
	.A(\eth_udp_inst|ip_send_inst|Add13~8_combout ),
	.B(\eth_udp_inst|ip_send_inst|LessThan1~3_combout ),
	.C(\eth_udp_inst|ip_send_inst|data_len [10]),
	.D(\eth_udp_inst|ip_send_inst|Add13~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .mask = 16'h8A08;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~5 (
	.A(\eth_udp_inst|ip_send_inst|LessThan1~2_combout ),
	.B(\eth_udp_inst|ip_send_inst|Add13~10_combout ),
	.C(\eth_udp_inst|ip_send_inst|LessThan1~4_combout ),
	.D(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~5_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .mask = 16'h7F01;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~6 (
	.A(\eth_udp_inst|ip_send_inst|Add13~16_combout ),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|LessThan1~5_combout ),
	.D(\eth_udp_inst|ip_send_inst|Add13~18_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~6_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .mask = 16'h0050;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~7 (
	.A(\eth_udp_inst|ip_send_inst|LessThan1~1_combout ),
	.B(\eth_udp_inst|ip_send_inst|LessThan1~6_combout ),
	.C(\eth_udp_inst|ip_send_inst|Add13~20_combout ),
	.D(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~7_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .mask = 16'h4544;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan2~0 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [13]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [11]),
	.C(\eth_udp_inst|ip_send_inst|data_cnt [12]),
	.D(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan2~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .mask = 16'h007F;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan2~1 (
	.A(\eth_udp_inst|ip_send_inst|Equal8~3_combout ),
	.B(\eth_udp_inst|ip_send_inst|data_len [10]),
	.C(\eth_udp_inst|ip_send_inst|data_cnt [8]),
	.D(\eth_udp_inst|ip_send_inst|data_cnt [9]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan2~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .mask = 16'h1333;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan2~2 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [8]),
	.B(\eth_udp_inst|ip_send_inst|Equal8~1_combout ),
	.C(\eth_udp_inst|ip_send_inst|Equal8~2_combout ),
	.D(\eth_udp_inst|ip_send_inst|data_cnt [9]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan2~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .mask = 16'h0015;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux13~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt [3]),
	.D(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux13~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .mask = 16'h1F00;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux13~1 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt [3]),
	.D(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux13~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .mask = 16'h2300;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux13~2 (
	.A(\eth_udp_inst|ip_send_inst|cnt [3]),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux13~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .mask = 16'h5500;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux13~3 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt [3]),
	.D(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux13~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .mask = 16'h1300;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux13~4 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt [3]),
	.D(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux13~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .mask = 16'h3700;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux16~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux16~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .mask = 16'h0008;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux17~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux17~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .mask = 16'h30BB;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux17~1 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Mux17~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux17~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .mask = 16'hC00C;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux20~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux20~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .mask = 16'h2E2C;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux21~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux21~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .mask = 16'h0F5D;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux24~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux24~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .mask = 16'hAF00;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux24~1 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|Mux24~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux24~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .mask = 16'h1A18;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux25~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux25~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .mask = 16'h1000;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux27~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux27~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .mask = 16'hFCF7;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux28~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux28~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .mask = 16'hF5A7;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux29~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux29~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .mask = 16'h0008;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux31~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux31~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .mask = 16'hFCF7;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux32~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|ip_udp_head[2][11]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux32~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .mask = 16'h0200;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux33~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[2][10]~q ),
	.D(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux33~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .mask = 16'hE200;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux35~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux35~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .mask = 16'h0CF0;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux35~1 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.D(\eth_udp_inst|ip_send_inst|Mux35~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux35~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .mask = 16'hBB98;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux36~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|ip_udp_head[2][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux36~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .mask = 16'h2420;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux37~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|ip_udp_head[2][14]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux37~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .mask = 16'hEDEF;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux39~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][12]~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|cnt [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux39~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .mask = 16'h0008;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux40~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[2][3]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux40~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .mask = 16'hC088;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux41~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|ip_udp_head[2][2]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux41~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .mask = 16'hC808;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux43~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][0]~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux43~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .mask = 16'hFDCF;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux44~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|ip_udp_head[2][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux44~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .mask = 16'h0400;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux45~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][6]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux45~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .mask = 16'h0400;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux47~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][4]~q ),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.D(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux47~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .mask = 16'hD800;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|always10~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always10~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|always10~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|always10~0 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|always10~0 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|always10~0 .mask = 16'h00C0;
defparam \eth_udp_inst|ip_send_inst|always10~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always10~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always10~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always10~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always10~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|always3~2 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always3~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|always3~2 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|always3~2 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|always3~2 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|always3~2 .mask = 16'h4040;
defparam \eth_udp_inst|ip_send_inst|always3~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|always3~3 (
	.A(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [4]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always3~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|always3~3 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|always3~3 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|always3~3 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|always3~3 .mask = 16'h0022;
defparam \eth_udp_inst|ip_send_inst|always3~3 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|always3~4 (
	.A(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.B(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always3~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|always3~4 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|always3~4 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|always3~4 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|always3~4 .mask = 16'h2222;
defparam \eth_udp_inst|ip_send_inst|always3~4 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|always7~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [3]),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always7~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|always7~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|always7~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|always7~0 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|always7~0 .mask = 16'h0040;
defparam \eth_udp_inst|ip_send_inst|always7~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|always7~1 (
	.A(\eth_udp_inst|ip_send_inst|always7~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|always10~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always7~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|always7~1 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|always7~1 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|always7~1 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|always7~1 .mask = 16'h0800;
defparam \eth_udp_inst|ip_send_inst|always7~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[0] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [16]),
	.B(\eth_udp_inst|ip_send_inst|check_sum [0]),
	.C(\eth_udp_inst|ip_send_inst|Add9~0_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [0]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y15_SIG ),
	.SyncReset(SyncReset_X28_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[0]~17_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[0]~18 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [0]));
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .mask = 16'h6688;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[10] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [10]),
	.C(\eth_udp_inst|ip_send_inst|Add9~20_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[9]~36 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [10]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y14_SIG ),
	.SyncReset(SyncReset_X28_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[10]~37_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[10]~38 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [10]));
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[11] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [11]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~22_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[10]~38 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [11]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y14_SIG ),
	.SyncReset(SyncReset_X28_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[11]~39_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[11]~40 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [11]));
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[12] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [12]),
	.C(\eth_udp_inst|ip_send_inst|Add9~24_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[11]~40 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [12]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y14_SIG ),
	.SyncReset(SyncReset_X28_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[12]~41_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[12]~42 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [12]));
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[13] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [13]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~26_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[12]~42 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [13]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y14_SIG ),
	.SyncReset(SyncReset_X28_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[13]~43_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[13]~44 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [13]));
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[14] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [14]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~28_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[13]~44 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [14]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y14_SIG ),
	.SyncReset(SyncReset_X28_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[14]~45_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[14]~46 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [14]));
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[15] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [15]),
	.C(\eth_udp_inst|ip_send_inst|Add9~30_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[14]~46 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [15]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y14_SIG ),
	.SyncReset(SyncReset_X28_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[15]~48_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[15]~49 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [15]));
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[16] (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~32_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[15]~49 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [16]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y14_SIG ),
	.SyncReset(SyncReset_X28_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[16]~52_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [16]));
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .mask = 16'h0F0F;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[17] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add9~34_combout ),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|Equal1~1_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [17]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum~51_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [17]));
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .mask = 16'hCC00;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[18] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Equal1~1_combout ),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|Add9~36_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [18]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum~50_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [18]));
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .mask = 16'hCC00;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[1] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [17]),
	.B(\eth_udp_inst|ip_send_inst|check_sum [1]),
	.C(\eth_udp_inst|ip_send_inst|Add9~2_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[0]~18 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [1]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y15_SIG ),
	.SyncReset(SyncReset_X28_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[1]~19_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[1]~20 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [1]));
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[2] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [2]),
	.B(\eth_udp_inst|ip_send_inst|check_sum [18]),
	.C(\eth_udp_inst|ip_send_inst|Add9~4_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[1]~20 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [2]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y15_SIG ),
	.SyncReset(SyncReset_X28_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[2]~21_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[2]~22 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [2]));
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[3] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [3]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~6_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[2]~22 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [3]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y15_SIG ),
	.SyncReset(SyncReset_X28_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[3]~23_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[3]~24 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [3]));
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[4] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [4]),
	.C(\eth_udp_inst|ip_send_inst|Add9~8_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[3]~24 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [4]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y15_SIG ),
	.SyncReset(SyncReset_X28_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[4]~25_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[4]~26 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [4]));
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[5] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [5]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~10_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[4]~26 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [5]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y15_SIG ),
	.SyncReset(SyncReset_X28_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[5]~27_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[5]~28 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [5]));
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[6] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [6]),
	.C(\eth_udp_inst|ip_send_inst|Add9~12_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[5]~28 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [6]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y15_SIG ),
	.SyncReset(SyncReset_X28_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[6]~29_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[6]~30 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [6]));
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[7] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [7]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~14_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[6]~30 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [7]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y15_SIG ),
	.SyncReset(SyncReset_X28_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[7]~31_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[7]~32 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [7]));
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[8] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [8]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~16_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[7]~32 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [8]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y14_SIG ),
	.SyncReset(SyncReset_X28_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[8]~33_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[8]~34 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [8]));
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[8]~47 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|always3~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[8]~47_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .mask = 16'h1500;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[9] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [9]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~18_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[8]~34 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [9]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y14_SIG ),
	.SyncReset(SyncReset_X28_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[9]~35_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[9]~36 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [9]));
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt[0] (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[3]~13_combout_X24_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|cnt[3]~11_combout__SyncReset_X24_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X24_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[0]~5_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt[0]~6 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt [0]));
defparam \eth_udp_inst|ip_send_inst|cnt[0] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .mask = 16'h55AA;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt[1] (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|cnt[0]~6 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[3]~13_combout_X24_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|cnt[3]~11_combout__SyncReset_X24_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X24_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[1]~7_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt[1]~8 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt [1]));
defparam \eth_udp_inst|ip_send_inst|cnt[1] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt[2] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|cnt[1]~8 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt [2]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[3]~13_combout_X24_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|cnt[3]~11_combout__SyncReset_X24_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X24_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[2]~9_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt[2]~10 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt [2]));
defparam \eth_udp_inst|ip_send_inst|cnt[2] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt[3] (
	.A(\eth_udp_inst|ip_send_inst|cnt [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|cnt[2]~10 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt [3]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[3]~13_combout_X24_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|cnt[3]~11_combout__SyncReset_X24_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X24_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[3]~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt[3]~15 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt [3]));
defparam \eth_udp_inst|ip_send_inst|cnt[3] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt[3]~11 (
	.A(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.B(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.C(\eth_udp_inst|ip_send_inst|always3~2_combout ),
	.D(\eth_udp_inst|ip_send_inst|always3~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[3]~11_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|cnt[3]~11 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~11 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~11 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~11 .mask = 16'hF444;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~11 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~11 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~11 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~11 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~11 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt[3]~12 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[3]~12_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|cnt[3]~12 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~12 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~12 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~12 .mask = 16'h7FFF;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~12 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~12 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt[3]~13 (
	.A(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt[3]~12_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[3]~13_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|cnt[3]~13 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~13 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~13 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~13 .mask = 16'hBABF;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~13 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~13 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~13 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~13 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3]~13 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt[4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt [4]),
	.Cin(\eth_udp_inst|ip_send_inst|cnt[3]~15 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt [4]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[3]~13_combout_X24_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|cnt[3]~11_combout__SyncReset_X24_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X24_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[4]~16_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|cnt [4]));
defparam \eth_udp_inst|ip_send_inst|cnt[4] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .mask = 16'hF00F;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_add[0] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt_add [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_add [0]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X22_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X22_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X22_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[0]~5_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt_add[0]~6 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt_add [0]));
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .mask = 16'h33CC;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt_add[1] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt_add [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|cnt_add[0]~6 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_add [1]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X22_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X22_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X22_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[1]~7_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt_add[1]~8 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt_add [1]));
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt_add[2] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt_add [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|cnt_add[1]~8 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_add [2]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X22_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X22_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X22_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[2]~9_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt_add[2]~10 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt_add [2]));
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt_add[3] (
	.A(\eth_udp_inst|ip_send_inst|cnt_add [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|cnt_add[2]~10 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_add [3]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X22_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X22_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X22_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[3]~11_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt_add[3]~12 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt_add [3]));
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt_add[4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt_add [4]),
	.Cin(\eth_udp_inst|ip_send_inst|cnt_add[3]~12 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_add [4]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X22_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X22_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X22_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[4]~13_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|cnt_add [4]));
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .mask = 16'hF00F;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_add[4]~15 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Equal8~6_combout ),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[4]~15_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .mask = 16'h00CC;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_send_bit[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout_X19_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X19_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_send_bit~5_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]));
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .mask = 16'h0F00;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_send_bit[1] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout_X19_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X19_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_send_bit~4_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]));
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .mask = 16'h3C00;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_send_bit[2] (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout_X19_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X19_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_send_bit~2_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]));
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .mask = 16'h7800;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 (
	.A(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .mask = 16'h0055;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.C(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .mask = 16'h72FA;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|crc_clr (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|send_end~q ),
	.D(\eth_udp_inst|ip_send_inst|crc_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Clk(\clk_25m~clkctrl_outclk_X22_Y19_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(SyncReset_X22_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X22_Y19_VCC),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data[28]~9_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|crc_clr~q ));
defparam \eth_udp_inst|ip_send_inst|crc_clr .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|crc_clr .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|crc_clr .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|crc_clr .mask = 16'hFFF0;
defparam \eth_udp_inst|ip_send_inst|crc_clr .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|crc_clr .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|crc_clr .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|crc_clr .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|crc_clr .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|crc_en (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|crc_en~q ),
	.Clk(\clk_25m~clkctrl_outclk_X23_Y18_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always13~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|crc_en~q ));
defparam \eth_udp_inst|ip_send_inst|crc_en .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|crc_en .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|crc_en .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|crc_en .mask = 16'hFFFC;
defparam \eth_udp_inst|ip_send_inst|crc_en .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|crc_en .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|crc_en .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|crc_en .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|crc_en .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[0] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [0]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[0]~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[0]~17 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [0]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .mask = 16'h55AA;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[10] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [10]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[9]~35 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [10]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[10]~36_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[10]~37 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [10]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[10]~41 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt[2]~40_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.C(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .mask = 16'h8088;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[11] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [11]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[10]~37 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [11]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[11]~42_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[11]~43 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [11]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[12] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [12]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[11]~43 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [12]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[12]~44_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[12]~45 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [12]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[13] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [13]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[12]~45 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [13]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[13]~46_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[13]~47 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [13]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[14] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [14]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[13]~47 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [14]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[14]~48_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[14]~49 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [14]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[15] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [15]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[14]~49 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [15]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[15]~50_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [15]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .mask = 16'h5A5A;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[1] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[0]~17 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [1]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[1]~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[1]~19 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [1]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[2] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[1]~19 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [2]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[2]~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[2]~21 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [2]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[2]~38 (
	.A(\eth_udp_inst|ip_send_inst|LessThan2~1_combout ),
	.B(\eth_udp_inst|ip_send_inst|Equal8~4_combout ),
	.C(\eth_udp_inst|ip_send_inst|LessThan2~2_combout ),
	.D(\eth_udp_inst|ip_send_inst|data_cnt [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[2]~38_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~38 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~38 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~38 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~38 .mask = 16'hC8CC;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~38 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~38 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~38 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~38 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~38 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[2]~39 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [15]),
	.B(\eth_udp_inst|ip_send_inst|LessThan2~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|data_len [10]),
	.D(\eth_udp_inst|ip_send_inst|data_cnt[2]~38_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[2]~39_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~39 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~39 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~39 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~39 .mask = 16'h5042;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~39 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~39 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~39 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~39 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~39 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[2]~40 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt[2]~39_combout ),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [14]),
	.C(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.D(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[2]~40_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~40 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~40 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~40 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~40 .mask = 16'hF2F7;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~40 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~40 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~40 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~40 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2]~40 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[3] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[2]~21 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [3]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[3]~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[3]~23 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [3]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[4] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[3]~23 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [4]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[4]~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[4]~25 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [4]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[5] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[4]~25 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [5]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[5]~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[5]~27 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [5]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[6] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[5]~27 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [6]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[6]~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[6]~29 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [6]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[7] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[6]~29 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [7]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[7]~30_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[7]~31 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [7]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[8] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [8]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[7]~31 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [8]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[8]~32_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[8]~33 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [8]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[9] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [9]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[8]~33 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [9]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X23_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[9]~34_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[9]~35 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [9]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_len[10] (
	.A(\LessThan0~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|send_en_r~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Clk(\clk_25m~clkctrl_outclk_X24_Y15_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|data_len[10]~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|data_len [10]));
defparam \eth_udp_inst|ip_send_inst|data_len[10] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .mask = 16'hF0F2;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data[0] (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~35_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~23_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~42_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.Clk(\clk_25m~clkctrl_outclk_X23_Y18_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~43_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|eth_tx_data [0]));
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .mask = 16'hFECC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data[1] (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~90_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~68_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.Clk(\clk_25m~clkctrl_outclk_X23_Y16_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~91_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|eth_tx_data [1]));
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .mask = 16'h0E02;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data[2] (
	.A(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~19_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.Clk(\clk_25m~clkctrl_outclk_X23_Y16_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~20_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|eth_tx_data [2]));
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .mask = 16'hFFA0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data[3] (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~65_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~64_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.Clk(\clk_25m~clkctrl_outclk_X23_Y16_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~66_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|eth_tx_data [3]));
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .mask = 16'hCCEC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~0 (
	.A(\eth_udp_inst|ip_send_inst|Mux13~1_combout ),
	.B(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|Mux13~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .mask = 16'hE3E0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~1 (
	.A(\eth_udp_inst|ip_send_inst|Mux13~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|Mux13~3_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .mask = 16'hCAF0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~10 (
	.A(\eth_udp_inst|crc32_inst|crc_data [21]),
	.B(\eth_udp_inst|crc32_inst|crc_data [17]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~9_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~10_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .mask = 16'hCAF0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~11 (
	.A(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~10_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~11_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .mask = 16'hA808;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~12 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~11_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.C(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.D(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~12_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .mask = 16'h00AE;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~13 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [15]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [13]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~13_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .mask = 16'hB9A8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~14 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [14]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~13_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [16]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~14_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .mask = 16'hEC2C;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~15 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [10]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [9]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~15_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .mask = 16'hD9C8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~16 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~15_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [11]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [12]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~16_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .mask = 16'hEA4A;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~17 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~14_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~16_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.D(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~17_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .mask = 16'hAC00;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~18 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~12_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~6_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~17_combout ),
	.D(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~18_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .mask = 16'hCCFE;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~19 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~1_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~18_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~19_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .mask = 16'h0B08;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~2 (
	.A(\eth_udp_inst|ip_send_inst|Mux33~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\eth_udp_inst|ip_send_inst|Mux41~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .mask = 16'hFC22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~21 (
	.A(\eth_udp_inst|ip_send_inst|cnt [3]),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~21_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .mask = 16'hC8EC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~22 (
	.A(\eth_udp_inst|ip_send_inst|cnt [3]),
	.B(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~21_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~22_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .mask = 16'h044C;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~23 (
	.A(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~22_combout ),
	.C(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~23_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .mask = 16'hA8A8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~24 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [14]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [13]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~24_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .mask = 16'hEE50;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~25 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~24_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [16]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [15]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~25_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .mask = 16'hE6C4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~26 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [10]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [9]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~26_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .mask = 16'hD9C8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~27 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [12]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~26_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [11]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~27_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .mask = 16'hBC8C;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~28 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~27_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~25_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~28_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .mask = 16'hC808;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~29 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|crc32_inst|crc_data [15]),
	.C(\eth_udp_inst|crc32_inst|crc_data [7]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~29_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .mask = 16'hAAE4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~3 (
	.A(\eth_udp_inst|ip_send_inst|Mux37~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|Mux45~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~2_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .mask = 16'hC5F0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~30 (
	.A(\eth_udp_inst|crc32_inst|crc_data [11]),
	.B(\eth_udp_inst|crc32_inst|crc_data [3]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~29_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~30_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .mask = 16'hCAF0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~31 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\eth_udp_inst|ip_send_inst|crc_en~q ),
	.D(\eth_udp_inst|crc32_inst|crc_data [27]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~31_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .mask = 16'hDD89;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~32 (
	.A(\eth_udp_inst|crc32_inst|crc_data [19]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.C(\eth_udp_inst|crc32_inst|crc_data [23]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~31_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~32_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .mask = 16'hBBC0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~33 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~32_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~30_combout ),
	.D(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~33_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .mask = 16'hE400;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~34 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.B(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~33_combout ),
	.D(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~34_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .mask = 16'h3032;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~35 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~28_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~34_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~35_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .mask = 16'h3330;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~36 (
	.A(\eth_udp_inst|ip_send_inst|Mux39~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.C(\eth_udp_inst|ip_send_inst|Mux35~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~36_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .mask = 16'hEE30;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~37 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~36_combout ),
	.B(\eth_udp_inst|ip_send_inst|Mux47~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|Mux43~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~37_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .mask = 16'h8DAA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~38 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~38_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .mask = 16'hDFF0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~39 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~39_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .mask = 16'hC500;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~4 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(\eth_udp_inst|ip_send_inst|Mux21~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|Mux17~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .mask = 16'hAAD8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~40 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~39_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~38_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~40_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .mask = 16'h88A9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~41 (
	.A(\eth_udp_inst|ip_send_inst|Mux27~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~40_combout ),
	.D(\eth_udp_inst|ip_send_inst|Mux31~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~41_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .mask = 16'h34F4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~42 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~41_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~37_combout ),
	.C(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~42_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .mask = 16'hC0A0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~44 (
	.A(\eth_udp_inst|ip_send_inst|cnt [3]),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~44_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .mask = 16'h5111;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~45 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~45_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .mask = 16'h0622;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~46 (
	.A(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.B(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~45_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~44_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~46_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .mask = 16'h8880;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~47 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|Mux40~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.D(\eth_udp_inst|ip_send_inst|Mux32~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~47_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .mask = 16'hADA8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~48 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~47_combout ),
	.B(\eth_udp_inst|ip_send_inst|Mux44~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.D(\eth_udp_inst|ip_send_inst|Mux36~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~48_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .mask = 16'hDA8A;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~49 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|Mux16~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|Mux20~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~49_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .mask = 16'hFA44;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~5 (
	.A(\eth_udp_inst|ip_send_inst|Mux25~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~4_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|Mux29~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~5_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .mask = 16'hEC2C;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~50 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|Mux28~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|Mux24~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~49_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~50_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .mask = 16'h77A0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~51 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~50_combout ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~48_combout ),
	.D(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~51_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .mask = 16'hE200;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~52 (
	.A(\eth_udp_inst|crc32_inst|crc_data [12]),
	.B(\eth_udp_inst|crc32_inst|crc_data [4]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~52_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .mask = 16'hF0CA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~53 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(\eth_udp_inst|crc32_inst|crc_data [8]),
	.C(\eth_udp_inst|crc32_inst|crc_data [0]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~52_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~53_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .mask = 16'hF588;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~54 (
	.A(\eth_udp_inst|crc32_inst|crc_data [24]),
	.B(\eth_udp_inst|crc32_inst|crc_next[28]~1_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~54_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .mask = 16'hFA03;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~55 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|crc32_inst|crc_data [16]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~54_combout ),
	.D(\eth_udp_inst|crc32_inst|crc_data [20]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~55_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .mask = 16'hDAD0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~56 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~55_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~53_combout ),
	.D(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~56_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .mask = 16'hE400;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~57 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~56_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.D(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~57_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .mask = 16'h00BA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~58 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [13]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [15]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~58_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .mask = 16'hAAE4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~59 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [16]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [14]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~58_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~59_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .mask = 16'hBBC0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~6 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~3_combout ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.C(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~6_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .mask = 16'hB080;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~60 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [10]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [9]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~60_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .mask = 16'hD9C8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~61 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [11]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a3__DataOutB [12]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~60_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~61_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .mask = 16'hF588;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~62 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.B(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~59_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~61_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~62_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .mask = 16'hC480;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~63 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~51_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~57_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~62_combout ),
	.D(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~63_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .mask = 16'hAAFE;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~65 (
	.A(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.B(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~65_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .mask = 16'h8000;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~67 (
	.A(\eth_udp_inst|ip_send_inst|Mux13~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|Mux13~3_combout ),
	.C(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~67_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .mask = 16'hFC0A;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~68 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~67_combout ),
	.B(\eth_udp_inst|ip_send_inst|Mux13~4_combout ),
	.C(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|Mux13~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~68_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .mask = 16'hDA8A;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~69 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][5]~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[2][13]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~69_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .mask = 16'hBBC0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~7 (
	.A(\eth_udp_inst|crc32_inst|crc_data [5]),
	.B(\eth_udp_inst|crc32_inst|crc_data [13]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~7_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .mask = 16'hF0AC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~70 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][9]~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~69_combout ),
	.D(\eth_udp_inst|ip_send_inst|ip_udp_head[2][1]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~70_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .mask = 16'hF2C2;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~71 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~70_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~71_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .mask = 16'h5CFA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~72 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~71_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~72_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .mask = 16'h0C30;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~73 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~q ),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~73_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .mask = 16'hAACC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~74 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~74_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .mask = 16'hBA00;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~75 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~75_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .mask = 16'h67CC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~76 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~75_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~76_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .mask = 16'h0DA0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~77 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~74_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~76_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~73_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~75_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~77_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .mask = 16'h88C8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~78 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~77_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~72_combout ),
	.D(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~78_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .mask = 16'hE400;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~79 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [15]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [13]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~79_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .mask = 16'hE3E0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~8 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~7_combout ),
	.B(\eth_udp_inst|crc32_inst|crc_data [9]),
	.C(\eth_udp_inst|crc32_inst|crc_data [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~8_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .mask = 16'hE4AA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~80 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [16]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [14]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~79_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~80_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .mask = 16'hBBC0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~81 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [9]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [10]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~81_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .mask = 16'hFC0A;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~82 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [11]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~81_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [12]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~82_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .mask = 16'hF858;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~83 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~82_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~80_combout ),
	.D(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~83_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .mask = 16'hE400;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~84 (
	.A(\eth_udp_inst|crc32_inst|crc_data [14]),
	.B(\eth_udp_inst|crc32_inst|crc_data [6]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~84_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .mask = 16'hF0CA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~85 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(\eth_udp_inst|crc32_inst|crc_data [10]),
	.C(\eth_udp_inst|crc32_inst|crc_data [2]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~84_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~85_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .mask = 16'hF588;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~86 (
	.A(\eth_udp_inst|crc32_inst|crc_data [26]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.D(\eth_udp_inst|ip_send_inst|crc_en~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~86_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .mask = 16'hE2E3;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~87 (
	.A(\eth_udp_inst|crc32_inst|crc_data [18]),
	.B(\eth_udp_inst|crc32_inst|crc_data [22]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~86_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~87_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .mask = 16'hAFC0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~88 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~87_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~85_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.D(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~88_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .mask = 16'hCA00;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~89 (
	.A(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.B(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~88_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~89_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .mask = 16'h3130;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~9 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\eth_udp_inst|crc32_inst|crc_next[29]~0_combout ),
	.D(\eth_udp_inst|crc32_inst|crc_data [25]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~9_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .mask = 16'hCD89;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~90 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~83_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~78_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~89_combout ),
	.D(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~90_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .mask = 16'hCCFE;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_en (
	.A(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|eth_tx_en~q ),
	.Clk(\clk_25m~clkctrl_outclk_X25_Y16_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always11~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|eth_tx_en~q ));
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .mask = 16'h5500;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] (
	.A(\eth_udp_inst|ip_send_inst|data_len [10]),
	.B(\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|always3~4_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.Clk(\clk_25m~clkctrl_outclk_X24_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X24_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~18_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .mask = 16'hE2F0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] (
	.A(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.B(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~q ),
	.Clk(\clk_25m~clkctrl_outclk_X24_Y15_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~53_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .mask = 16'hD2D2;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~21_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~22 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .mask = 16'h6688;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~22 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~23_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~24 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~24 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~25_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~26 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~26 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~27_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~28 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~28 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~29_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~30 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~30 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~31_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~32 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~32 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~33_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~34 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~34 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~35_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~36 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~36 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~37_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~38 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~38 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~39_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~40 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~40 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~41_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~42 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~42 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~43_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~44 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~44 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~45_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~46 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~46 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~47_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~48 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~q ),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~48 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X25_Y17_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~58_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .mask = 16'hF00F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [0]),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][0]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~49_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][0]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .mask = 16'h3033;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] (
	.A(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.B(\eth_udp_inst|ip_send_inst|check_sum [10]),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][10]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~19_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][10]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .mask = 16'h3131;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [11]),
	.B(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][11]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~56_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][11]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .mask = 16'h5151;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] (
	.A(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.B(\eth_udp_inst|ip_send_inst|check_sum [12]),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][12]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~50_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][12]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .mask = 16'h3131;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [13]),
	.B(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][13]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~62_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][13]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .mask = 16'h5151;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [14]),
	.B(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][14]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~15_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][14]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .mask = 16'h5151;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.C(\eth_udp_inst|ip_send_inst|check_sum [15]),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][15]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~54_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][15]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .mask = 16'h0C0F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [1]),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][1]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~60_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][1]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .mask = 16'h3033;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.C(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.D(\eth_udp_inst|ip_send_inst|check_sum [2]),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][2]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~17_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][2]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .mask = 16'h00CF;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [3]),
	.B(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][3]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~55_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][3]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .mask = 16'h5151;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [4]),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][4]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~52_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][4]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .mask = 16'h3033;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.C(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.D(\eth_udp_inst|ip_send_inst|check_sum [5]),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][5]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~63_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][5]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .mask = 16'h00CF;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [6]),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][6]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~20_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][6]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .mask = 16'h3033;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [7]),
	.B(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][7]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~57_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][7]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .mask = 16'h4455;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [8]),
	.B(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~51_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .mask = 16'h5151;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 (
	.A(\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.B(\eth_udp_inst|ip_send_inst|always3~3_combout ),
	.C(\eth_udp_inst|ip_send_inst|always3~2_combout ),
	.D(\eth_udp_inst|ip_send_inst|always3~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .mask = 16'h5540;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [9]),
	.B(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][9]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X28_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X28_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~61_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][9]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .mask = 16'h5151;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|packet_head[7][7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.Clk(\clk_25m~clkctrl_outclk_X23_Y16_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|packet_head[7][7]~feeder_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ));
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .mask = 16'hFFFF;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|read_data_req (
	.A(\eth_udp_inst|ip_send_inst|always10~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|Equal8~6_combout ),
	.C(\eth_udp_inst|ip_send_inst|always7~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|read_data_req~q ),
	.Clk(\clk_25m~clkctrl_outclk_X23_Y18_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|read_data_req~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|read_data_req~q ));
defparam \eth_udp_inst|ip_send_inst|read_data_req .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|read_data_req .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|read_data_req .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|read_data_req .mask = 16'hF2F0;
defparam \eth_udp_inst|ip_send_inst|read_data_req .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|read_data_req .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|read_data_req .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|read_data_req .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|read_data_req .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|send_en_r (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|send_en_r~q ),
	.Clk(\clk_25m~clkctrl_outclk_X24_Y15_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\LessThan0~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|send_en_r~q ));
defparam \eth_udp_inst|ip_send_inst|send_en_r .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|send_en_r .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|send_en_r .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|send_en_r .mask = 16'hFAF8;
defparam \eth_udp_inst|ip_send_inst|send_en_r .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_en_r .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_en_r .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_en_r .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_en_r .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|send_end (
	.A(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|send_end~q ),
	.Clk(\clk_25m~clkctrl_outclk_X23_Y18_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always16~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|send_end~q ));
defparam \eth_udp_inst|ip_send_inst|send_end .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|send_end .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|send_end .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|send_end .mask = 16'h8000;
defparam \eth_udp_inst|ip_send_inst|send_end .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_end .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_end .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_end .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_end .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.CHECK_SUM (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X25_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ));
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .mask = 16'h00FF;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.CRC (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y18_SIG ),
	.SyncReset(SyncReset_X23_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y18_VCC),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~5_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.CRC~q ));
defparam \eth_udp_inst|ip_send_inst|state.CRC .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|state.CRC .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|state.CRC .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|state.CRC .mask = 16'hA000;
defparam \eth_udp_inst|ip_send_inst|state.CRC .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.CRC .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.CRC .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.CRC .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.CRC .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.ETH_HEAD (
	.A(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~46_combout ),
	.C(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~63_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(SyncReset_X23_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y16_VCC),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~64_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ));
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .mask = 16'h4544;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.IDLE (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X24_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|state.IDLE~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.IDLE~q ));
defparam \eth_udp_inst|ip_send_inst|state.IDLE .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .mask = 16'h0F0F;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD (
	.A(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.B(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.C(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y18_SIG ),
	.SyncReset(SyncReset_X23_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y18_VCC),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ));
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .mask = 16'hFEFF;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.PACKET_HEAD (
	.A(\eth_udp_inst|ip_send_inst|cnt [3]),
	.B(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(SyncReset_X23_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y16_VCC),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~1_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ));
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .mask = 16'h5088;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.SEND_DATA (
	.A(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.B(\eth_udp_inst|ip_send_inst|LessThan1~7_combout ),
	.C(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_add[4]~15_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y18_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y18_SIG ),
	.SyncReset(SyncReset_X23_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y18_VCC),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ));
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .mask = 16'hE0A0;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|sw_en (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\eth_udp_inst|ip_send_inst|sw_en~6_combout ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~4_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Clk(\clk_25m~clkctrl_outclk_X24_Y15_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~7_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|sw_en~q ));
defparam \eth_udp_inst|ip_send_inst|sw_en .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|sw_en .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|sw_en .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|sw_en .mask = 16'hFF30;
defparam \eth_udp_inst|ip_send_inst|sw_en .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|sw_en~0 (
	.A(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .mask = 16'h0080;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|sw_en~2 (
	.A(\eth_udp_inst|ip_send_inst|sw_en~1_combout ),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .mask = 16'h8000;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|sw_en~3 (
	.A(\eth_udp_inst|ip_send_inst|cnt [4]),
	.B(\eth_udp_inst|ip_send_inst|sw_en~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|always7~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .mask = 16'hF5F4;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|sw_en~4 (
	.A(\LessThan0~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.C(\eth_udp_inst|ip_send_inst|sw_en~3_combout ),
	.D(\eth_udp_inst|ip_send_inst|send_en_r~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .mask = 16'hF0F2;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|sw_en~6 (
	.A(\eth_udp_inst|ip_send_inst|sw_en~5_combout ),
	.B(\eth_udp_inst|ip_send_inst|Equal8~6_combout ),
	.C(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.D(\eth_udp_inst|ip_send_inst|LessThan1~7_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~6_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .mask = 16'hAAEA;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .CarryEnb = 1'b1;

alta_slice led_r(
	.A(\Equal0~4_combout ),
	.B(\Equal0~5_combout ),
	.C(vcc),
	.D(\Equal0~7_combout ),
	.Cin(),
	.Qin(\led_r~q ),
	.Clk(\clk~inputclkctrl_outclk_X11_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\led_r~0_combout ),
	.Cout(),
	.Q(\led_r~q ));
defparam led_r.coord_x = 1;
defparam led_r.coord_y = 9;
defparam led_r.coord_z = 6;
defparam led_r.mask = 16'h78F0;
defparam led_r.modeMux = 1'b0;
defparam led_r.FeedbackMux = 1'b1;
defparam led_r.ShiftMux = 1'b0;
defparam led_r.BypassEn = 1'b0;
defparam led_r.CarryEnb = 1'b1;

alta_dio \led~output (
	.padio(led),
	.datain(\led_r~q ),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \led~output .coord_x = 0;
defparam \led~output .coord_y = 15;
defparam \led~output .coord_z = 2;
defparam \led~output .IN_ASYNC_MODE = 1'b0;
defparam \led~output .IN_SYNC_MODE = 1'b0;
defparam \led~output .IN_POWERUP = 1'b0;
defparam \led~output .IN_ASYNC_DISABLE = 1'b0;
defparam \led~output .IN_SYNC_DISABLE = 1'b0;
defparam \led~output .OUT_REG_MODE = 1'b0;
defparam \led~output .OUT_ASYNC_MODE = 1'b0;
defparam \led~output .OUT_SYNC_MODE = 1'b0;
defparam \led~output .OUT_POWERUP = 1'b0;
defparam \led~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \led~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \led~output .OUT_SYNC_DISABLE = 1'b0;
defparam \led~output .OUT_DDIO = 1'b0;
defparam \led~output .OE_REG_MODE = 1'b0;
defparam \led~output .OE_ASYNC_MODE = 1'b0;
defparam \led~output .OE_SYNC_MODE = 1'b0;
defparam \led~output .OE_POWERUP = 1'b0;
defparam \led~output .OE_CLKEN_DISABLE = 1'b0;
defparam \led~output .OE_ASYNC_DISABLE = 1'b0;
defparam \led~output .OE_SYNC_DISABLE = 1'b0;
defparam \led~output .OE_DDIO = 1'b0;
defparam \led~output .CFG_TRI_INPUT = 1'b0;
defparam \led~output .CFG_PULL_UP = 1'b0;
defparam \led~output .CFG_OPEN_DRAIN = 1'b0;
defparam \led~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \led~output .CFG_PDRV = 7'b0011010;
defparam \led~output .CFG_NDRV = 7'b0011000;
defparam \led~output .CFG_KEEP = 2'b00;
defparam \led~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \led~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \led~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \led~output .CFG_LVDS_IN_EN = 1'b0;
defparam \led~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \led~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \led~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \led~output .CFG_OSCDIV = 2'b00;
defparam \led~output .CFG_ROCTUSR = 1'b0;
defparam \led~output .CFG_SEL_CUA = 1'b0;
defparam \led~output .CFG_ROCT_EN = 1'b0;
defparam \led~output .INPUT_ONLY = 1'b0;
defparam \led~output .DPCLK_DELAY = 4'b0000;
defparam \led~output .OUT_DELAY = 1'b0;
defparam \led~output .IN_DATA_DELAY = 3'b000;
defparam \led~output .IN_REG_DELAY = 3'b000;

alta_slice \mii_to_rmii_inst|eth_tx_data[0] (
	.A(\mii_to_rmii_inst|eth_tx_data_reg [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\mii_to_rmii_inst|eth_tx_data [0]),
	.Clk(\e_rxclk~input_o_X23_Y19_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|eth_tx_data[0]~feeder_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|eth_tx_data [0]));
defparam \mii_to_rmii_inst|eth_tx_data[0] .coord_x = 21;
defparam \mii_to_rmii_inst|eth_tx_data[0] .coord_y = 17;
defparam \mii_to_rmii_inst|eth_tx_data[0] .coord_z = 12;
defparam \mii_to_rmii_inst|eth_tx_data[0] .mask = 16'hAAAA;
defparam \mii_to_rmii_inst|eth_tx_data[0] .modeMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[0] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[0] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[0] .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[0] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|eth_tx_data[1] (
	.A(),
	.B(),
	.C(\mii_to_rmii_inst|eth_tx_data_reg [1]),
	.D(),
	.Cin(),
	.Qin(\mii_to_rmii_inst|eth_tx_data [1]),
	.Clk(\e_rxclk~input_o_X23_Y19_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(SyncReset_X23_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y19_VCC),
	.LutOut(),
	.Cout(),
	.Q(\mii_to_rmii_inst|eth_tx_data [1]));
defparam \mii_to_rmii_inst|eth_tx_data[1] .coord_x = 21;
defparam \mii_to_rmii_inst|eth_tx_data[1] .coord_y = 17;
defparam \mii_to_rmii_inst|eth_tx_data[1] .coord_z = 13;
defparam \mii_to_rmii_inst|eth_tx_data[1] .mask = 16'hFFFF;
defparam \mii_to_rmii_inst|eth_tx_data[1] .modeMux = 1'b1;
defparam \mii_to_rmii_inst|eth_tx_data[1] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[1] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[1] .BypassEn = 1'b1;
defparam \mii_to_rmii_inst|eth_tx_data[1] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|eth_tx_data_reg[0] (
	.A(\mii_to_rmii_inst|rd_flag~q ),
	.B(\mii_to_rmii_inst|tx_data_reg [0]),
	.C(vcc),
	.D(\mii_to_rmii_inst|tx_data_reg [2]),
	.Cin(),
	.Qin(\mii_to_rmii_inst|eth_tx_data_reg [0]),
	.Clk(\e_rxclk~input_o__mii_to_rmii_inst|tx_dv_reg~q_X23_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|eth_tx_data_reg~0_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|eth_tx_data_reg [0]));
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .coord_x = 21;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .coord_y = 17;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .coord_z = 3;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .mask = 16'hEE44;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .modeMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|eth_tx_data_reg[1] (
	.A(\mii_to_rmii_inst|rd_flag~q ),
	.B(\mii_to_rmii_inst|tx_data_reg [1]),
	.C(\mii_to_rmii_inst|tx_data_reg [3]),
	.D(vcc),
	.Cin(),
	.Qin(\mii_to_rmii_inst|eth_tx_data_reg [1]),
	.Clk(\e_rxclk~input_o__mii_to_rmii_inst|tx_dv_reg~q_X23_Y19_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|eth_tx_data_reg~1_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|eth_tx_data_reg [1]));
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .coord_x = 21;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .coord_y = 17;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .coord_z = 11;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .mask = 16'hE4E4;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .modeMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|eth_tx_dv (
	.A(vcc),
	.B(\mii_to_rmii_inst|tx_dv_reg~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\mii_to_rmii_inst|eth_tx_dv~q ),
	.Clk(\e_rxclk~input_o_X23_Y19_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|eth_tx_dv~feeder_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|eth_tx_dv~q ));
defparam \mii_to_rmii_inst|eth_tx_dv .coord_x = 21;
defparam \mii_to_rmii_inst|eth_tx_dv .coord_y = 17;
defparam \mii_to_rmii_inst|eth_tx_dv .coord_z = 0;
defparam \mii_to_rmii_inst|eth_tx_dv .mask = 16'hCCCC;
defparam \mii_to_rmii_inst|eth_tx_dv .modeMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_dv .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_dv .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_dv .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_dv .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|rd_flag (
	.A(vcc),
	.B(\mii_to_rmii_inst|tx_dv_reg~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\mii_to_rmii_inst|rd_flag~q ),
	.Clk(\e_rxclk~input_o_X23_Y19_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|rd_flag~0_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|rd_flag~q ));
defparam \mii_to_rmii_inst|rd_flag .coord_x = 21;
defparam \mii_to_rmii_inst|rd_flag .coord_y = 17;
defparam \mii_to_rmii_inst|rd_flag .coord_z = 15;
defparam \mii_to_rmii_inst|rd_flag .mask = 16'h0C0C;
defparam \mii_to_rmii_inst|rd_flag .modeMux = 1'b0;
defparam \mii_to_rmii_inst|rd_flag .FeedbackMux = 1'b1;
defparam \mii_to_rmii_inst|rd_flag .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|rd_flag .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|rd_flag .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|tx_data_reg[0] (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.D(vcc),
	.Cin(),
	.Qin(\mii_to_rmii_inst|tx_data_reg [0]),
	.Clk(\e_rxclk~input_o_X23_Y19_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|tx_data_reg[0]~feeder_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|tx_data_reg [0]));
defparam \mii_to_rmii_inst|tx_data_reg[0] .coord_x = 21;
defparam \mii_to_rmii_inst|tx_data_reg[0] .coord_y = 17;
defparam \mii_to_rmii_inst|tx_data_reg[0] .coord_z = 14;
defparam \mii_to_rmii_inst|tx_data_reg[0] .mask = 16'hF0F0;
defparam \mii_to_rmii_inst|tx_data_reg[0] .modeMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[0] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[0] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[0] .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[0] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|tx_data_reg[1] (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.D(vcc),
	.Cin(),
	.Qin(\mii_to_rmii_inst|tx_data_reg [1]),
	.Clk(\e_rxclk~input_o_X23_Y19_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|tx_data_reg[1]~feeder_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|tx_data_reg [1]));
defparam \mii_to_rmii_inst|tx_data_reg[1] .coord_x = 21;
defparam \mii_to_rmii_inst|tx_data_reg[1] .coord_y = 17;
defparam \mii_to_rmii_inst|tx_data_reg[1] .coord_z = 4;
defparam \mii_to_rmii_inst|tx_data_reg[1] .mask = 16'hF0F0;
defparam \mii_to_rmii_inst|tx_data_reg[1] .modeMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[1] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[1] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[1] .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[1] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|tx_data_reg[2] (
	.A(),
	.B(),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.D(),
	.Cin(),
	.Qin(\mii_to_rmii_inst|tx_data_reg [2]),
	.Clk(\e_rxclk~input_o_X23_Y19_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(SyncReset_X23_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y19_VCC),
	.LutOut(),
	.Cout(),
	.Q(\mii_to_rmii_inst|tx_data_reg [2]));
defparam \mii_to_rmii_inst|tx_data_reg[2] .coord_x = 21;
defparam \mii_to_rmii_inst|tx_data_reg[2] .coord_y = 17;
defparam \mii_to_rmii_inst|tx_data_reg[2] .coord_z = 8;
defparam \mii_to_rmii_inst|tx_data_reg[2] .mask = 16'hFFFF;
defparam \mii_to_rmii_inst|tx_data_reg[2] .modeMux = 1'b1;
defparam \mii_to_rmii_inst|tx_data_reg[2] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[2] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[2] .BypassEn = 1'b1;
defparam \mii_to_rmii_inst|tx_data_reg[2] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|tx_data_reg[3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.Cin(),
	.Qin(\mii_to_rmii_inst|tx_data_reg [3]),
	.Clk(\e_rxclk~input_o_X23_Y19_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|tx_data_reg[3]~feeder_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|tx_data_reg [3]));
defparam \mii_to_rmii_inst|tx_data_reg[3] .coord_x = 21;
defparam \mii_to_rmii_inst|tx_data_reg[3] .coord_y = 17;
defparam \mii_to_rmii_inst|tx_data_reg[3] .coord_z = 1;
defparam \mii_to_rmii_inst|tx_data_reg[3] .mask = 16'hFF00;
defparam \mii_to_rmii_inst|tx_data_reg[3] .modeMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[3] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[3] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[3] .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[3] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|tx_dv_reg (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_en~q ),
	.D(vcc),
	.Cin(),
	.Qin(\mii_to_rmii_inst|tx_dv_reg~q ),
	.Clk(\e_rxclk~input_o_X23_Y19_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|tx_dv_reg~feeder_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|tx_dv_reg~q ));
defparam \mii_to_rmii_inst|tx_dv_reg .coord_x = 21;
defparam \mii_to_rmii_inst|tx_dv_reg .coord_y = 17;
defparam \mii_to_rmii_inst|tx_dv_reg .coord_z = 7;
defparam \mii_to_rmii_inst|tx_dv_reg .mask = 16'hF0F0;
defparam \mii_to_rmii_inst|tx_dv_reg .modeMux = 1'b0;
defparam \mii_to_rmii_inst|tx_dv_reg .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|tx_dv_reg .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|tx_dv_reg .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|tx_dv_reg .CarryEnb = 1'b1;

alta_slice \reset_init[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(reset_init[0]),
	.Clk(\clk~inputclkctrl_outclk__reset_init[5]_X12_Y12_SIG_INV ),
	.AsyncReset(AsyncReset_X12_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\reset_init[0]~1_combout ),
	.Cout(),
	.Q(reset_init[0]));
defparam \reset_init[0] .coord_x = 47;
defparam \reset_init[0] .coord_y = 15;
defparam \reset_init[0] .coord_z = 5;
defparam \reset_init[0] .mask = 16'h0F0F;
defparam \reset_init[0] .modeMux = 1'b0;
defparam \reset_init[0] .FeedbackMux = 1'b1;
defparam \reset_init[0] .ShiftMux = 1'b0;
defparam \reset_init[0] .BypassEn = 1'b0;
defparam \reset_init[0] .CarryEnb = 1'b1;

alta_slice \reset_init[1] (
	.A(reset_init[0]),
	.B(reset_init[1]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(reset_init[1]),
	.Clk(\clk~inputclkctrl_outclk__reset_init[5]_X12_Y12_SIG_INV ),
	.AsyncReset(AsyncReset_X12_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Add0~0_combout ),
	.Cout(\Add0~1 ),
	.Q(reset_init[1]));
defparam \reset_init[1] .coord_x = 47;
defparam \reset_init[1] .coord_y = 15;
defparam \reset_init[1] .coord_z = 8;
defparam \reset_init[1] .mask = 16'h6688;
defparam \reset_init[1] .modeMux = 1'b0;
defparam \reset_init[1] .FeedbackMux = 1'b0;
defparam \reset_init[1] .ShiftMux = 1'b0;
defparam \reset_init[1] .BypassEn = 1'b0;
defparam \reset_init[1] .CarryEnb = 1'b0;

alta_slice \reset_init[2] (
	.A(vcc),
	.B(reset_init[2]),
	.C(vcc),
	.D(vcc),
	.Cin(\Add0~1 ),
	.Qin(reset_init[2]),
	.Clk(\clk~inputclkctrl_outclk__reset_init[5]_X12_Y12_SIG_INV ),
	.AsyncReset(AsyncReset_X12_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Add0~2_combout ),
	.Cout(\Add0~3 ),
	.Q(reset_init[2]));
defparam \reset_init[2] .coord_x = 47;
defparam \reset_init[2] .coord_y = 15;
defparam \reset_init[2] .coord_z = 9;
defparam \reset_init[2] .mask = 16'h3C3F;
defparam \reset_init[2] .modeMux = 1'b1;
defparam \reset_init[2] .FeedbackMux = 1'b0;
defparam \reset_init[2] .ShiftMux = 1'b0;
defparam \reset_init[2] .BypassEn = 1'b0;
defparam \reset_init[2] .CarryEnb = 1'b0;

alta_slice \reset_init[3] (
	.A(vcc),
	.B(reset_init[3]),
	.C(vcc),
	.D(vcc),
	.Cin(\Add0~3 ),
	.Qin(reset_init[3]),
	.Clk(\clk~inputclkctrl_outclk__reset_init[5]_X12_Y12_SIG_INV ),
	.AsyncReset(AsyncReset_X12_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Add0~4_combout ),
	.Cout(\Add0~5 ),
	.Q(reset_init[3]));
defparam \reset_init[3] .coord_x = 47;
defparam \reset_init[3] .coord_y = 15;
defparam \reset_init[3] .coord_z = 10;
defparam \reset_init[3] .mask = 16'hC30C;
defparam \reset_init[3] .modeMux = 1'b1;
defparam \reset_init[3] .FeedbackMux = 1'b0;
defparam \reset_init[3] .ShiftMux = 1'b0;
defparam \reset_init[3] .BypassEn = 1'b0;
defparam \reset_init[3] .CarryEnb = 1'b0;

alta_slice \reset_init[4] (
	.A(reset_init[4]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\Add0~5 ),
	.Qin(reset_init[4]),
	.Clk(\clk~inputclkctrl_outclk__reset_init[5]_X12_Y12_SIG_INV ),
	.AsyncReset(AsyncReset_X12_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Add0~6_combout ),
	.Cout(\Add0~7 ),
	.Q(reset_init[4]));
defparam \reset_init[4] .coord_x = 47;
defparam \reset_init[4] .coord_y = 15;
defparam \reset_init[4] .coord_z = 11;
defparam \reset_init[4] .mask = 16'h5A5F;
defparam \reset_init[4] .modeMux = 1'b1;
defparam \reset_init[4] .FeedbackMux = 1'b0;
defparam \reset_init[4] .ShiftMux = 1'b0;
defparam \reset_init[4] .BypassEn = 1'b0;
defparam \reset_init[4] .CarryEnb = 1'b0;

alta_slice \reset_init[5] (
	.A(vcc),
	.B(\Add0~8_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(reset_init[5]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y12_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\reset_init[5]~0_combout ),
	.Cout(),
	.Q(reset_init[5]));
defparam \reset_init[5] .coord_x = 47;
defparam \reset_init[5] .coord_y = 15;
defparam \reset_init[5] .coord_z = 4;
defparam \reset_init[5] .mask = 16'hFCFC;
defparam \reset_init[5] .modeMux = 1'b0;
defparam \reset_init[5] .FeedbackMux = 1'b1;
defparam \reset_init[5] .ShiftMux = 1'b0;
defparam \reset_init[5] .BypassEn = 1'b0;
defparam \reset_init[5] .CarryEnb = 1'b1;

alta_io_gclk \reset_init[5]~clkctrl (
	.inclk(reset_init[5]),
	.outclk(\reset_init[5]~clkctrl_outclk ));
defparam \reset_init[5]~clkctrl .coord_x = 49;
defparam \reset_init[5]~clkctrl .coord_y = 15;
defparam \reset_init[5]~clkctrl .coord_z = 3;

alta_dio \rst_n~input (
	.padio(rst_n),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\rst_n~input_o ),
	.regout());
defparam \rst_n~input .coord_x = 49;
defparam \rst_n~input .coord_y = 15;
defparam \rst_n~input .coord_z = 0;
defparam \rst_n~input .IN_ASYNC_MODE = 1'b0;
defparam \rst_n~input .IN_SYNC_MODE = 1'b0;
defparam \rst_n~input .IN_POWERUP = 1'b0;
defparam \rst_n~input .IN_ASYNC_DISABLE = 1'b0;
defparam \rst_n~input .IN_SYNC_DISABLE = 1'b0;
defparam \rst_n~input .OUT_REG_MODE = 1'b0;
defparam \rst_n~input .OUT_ASYNC_MODE = 1'b0;
defparam \rst_n~input .OUT_SYNC_MODE = 1'b0;
defparam \rst_n~input .OUT_POWERUP = 1'b0;
defparam \rst_n~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \rst_n~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \rst_n~input .OUT_SYNC_DISABLE = 1'b0;
defparam \rst_n~input .OUT_DDIO = 1'b0;
defparam \rst_n~input .OE_REG_MODE = 1'b0;
defparam \rst_n~input .OE_ASYNC_MODE = 1'b0;
defparam \rst_n~input .OE_SYNC_MODE = 1'b0;
defparam \rst_n~input .OE_POWERUP = 1'b0;
defparam \rst_n~input .OE_CLKEN_DISABLE = 1'b0;
defparam \rst_n~input .OE_ASYNC_DISABLE = 1'b0;
defparam \rst_n~input .OE_SYNC_DISABLE = 1'b0;
defparam \rst_n~input .OE_DDIO = 1'b0;
defparam \rst_n~input .CFG_TRI_INPUT = 1'b0;
defparam \rst_n~input .CFG_PULL_UP = 1'b0;
defparam \rst_n~input .CFG_OPEN_DRAIN = 1'b0;
defparam \rst_n~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \rst_n~input .CFG_PDRV = 7'b0010000;
defparam \rst_n~input .CFG_NDRV = 7'b0010000;
defparam \rst_n~input .CFG_KEEP = 2'b00;
defparam \rst_n~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \rst_n~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \rst_n~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \rst_n~input .CFG_LVDS_IN_EN = 1'b0;
defparam \rst_n~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \rst_n~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \rst_n~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \rst_n~input .CFG_OSCDIV = 2'b00;
defparam \rst_n~input .CFG_ROCTUSR = 1'b0;
defparam \rst_n~input .CFG_SEL_CUA = 1'b0;
defparam \rst_n~input .CFG_ROCT_EN = 1'b0;
defparam \rst_n~input .INPUT_ONLY = 1'b1;
defparam \rst_n~input .DPCLK_DELAY = 4'b0000;
defparam \rst_n~input .OUT_DELAY = 1'b0;
defparam \rst_n~input .IN_DATA_DELAY = 3'b000;
defparam \rst_n~input .IN_REG_DELAY = 3'b000;

alta_syncctrl syncload_ctrl_X12_Y13(
	.Din(),
	.Dout(SyncLoad_X12_Y13_VCC));
defparam syncload_ctrl_X12_Y13.coord_x = 16;
defparam syncload_ctrl_X12_Y13.coord_y = 13;
defparam syncload_ctrl_X12_Y13.coord_z = 1;
defparam syncload_ctrl_X12_Y13.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X12_Y14(
	.Din(),
	.Dout(SyncLoad_X12_Y14_GND));
defparam syncload_ctrl_X12_Y14.coord_x = 2;
defparam syncload_ctrl_X12_Y14.coord_y = 9;
defparam syncload_ctrl_X12_Y14.coord_z = 1;
defparam syncload_ctrl_X12_Y14.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X12_Y15(
	.Din(),
	.Dout(SyncLoad_X12_Y15_GND));
defparam syncload_ctrl_X12_Y15.coord_x = 2;
defparam syncload_ctrl_X12_Y15.coord_y = 10;
defparam syncload_ctrl_X12_Y15.coord_z = 1;
defparam syncload_ctrl_X12_Y15.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X13_Y12(
	.Din(),
	.Dout(SyncLoad_X13_Y12_VCC));
defparam syncload_ctrl_X13_Y12.coord_x = 15;
defparam syncload_ctrl_X13_Y12.coord_y = 16;
defparam syncload_ctrl_X13_Y12.coord_z = 1;
defparam syncload_ctrl_X13_Y12.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X14_Y12(
	.Din(),
	.Dout(SyncLoad_X14_Y12_VCC));
defparam syncload_ctrl_X14_Y12.coord_x = 17;
defparam syncload_ctrl_X14_Y12.coord_y = 16;
defparam syncload_ctrl_X14_Y12.coord_z = 1;
defparam syncload_ctrl_X14_Y12.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X14_Y13(
	.Din(),
	.Dout(SyncLoad_X14_Y13_VCC));
defparam syncload_ctrl_X14_Y13.coord_x = 17;
defparam syncload_ctrl_X14_Y13.coord_y = 13;
defparam syncload_ctrl_X14_Y13.coord_z = 1;
defparam syncload_ctrl_X14_Y13.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X14_Y17(
	.Din(),
	.Dout(SyncLoad_X14_Y17_GND));
defparam syncload_ctrl_X14_Y17.coord_x = 10;
defparam syncload_ctrl_X14_Y17.coord_y = 15;
defparam syncload_ctrl_X14_Y17.coord_z = 1;
defparam syncload_ctrl_X14_Y17.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X16_Y11(
	.Din(),
	.Dout(SyncLoad_X16_Y11_VCC));
defparam syncload_ctrl_X16_Y11.coord_x = 17;
defparam syncload_ctrl_X16_Y11.coord_y = 15;
defparam syncload_ctrl_X16_Y11.coord_z = 1;
defparam syncload_ctrl_X16_Y11.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X16_Y12(
	.Din(),
	.Dout(SyncLoad_X16_Y12_VCC));
defparam syncload_ctrl_X16_Y12.coord_x = 16;
defparam syncload_ctrl_X16_Y12.coord_y = 16;
defparam syncload_ctrl_X16_Y12.coord_z = 1;
defparam syncload_ctrl_X16_Y12.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X16_Y13(
	.Din(),
	.Dout(SyncLoad_X16_Y13_VCC));
defparam syncload_ctrl_X16_Y13.coord_x = 17;
defparam syncload_ctrl_X16_Y13.coord_y = 14;
defparam syncload_ctrl_X16_Y13.coord_z = 1;
defparam syncload_ctrl_X16_Y13.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X17_Y13(
	.Din(),
	.Dout(SyncLoad_X17_Y13_VCC));
defparam syncload_ctrl_X17_Y13.coord_x = 16;
defparam syncload_ctrl_X17_Y13.coord_y = 15;
defparam syncload_ctrl_X17_Y13.coord_z = 1;
defparam syncload_ctrl_X17_Y13.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X1_Y17(
	.Din(),
	.Dout(SyncLoad_X1_Y17_GND));
defparam syncload_ctrl_X1_Y17.coord_x = 11;
defparam syncload_ctrl_X1_Y17.coord_y = 16;
defparam syncload_ctrl_X1_Y17.coord_z = 1;
defparam syncload_ctrl_X1_Y17.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X1_Y7(
	.Din(),
	.Dout(SyncLoad_X1_Y7_VCC));
defparam syncload_ctrl_X1_Y7.coord_x = 8;
defparam syncload_ctrl_X1_Y7.coord_y = 12;
defparam syncload_ctrl_X1_Y7.coord_z = 1;
defparam syncload_ctrl_X1_Y7.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X22_Y16(
	.Din(),
	.Dout(SyncLoad_X22_Y16_GND));
defparam syncload_ctrl_X22_Y16.coord_x = 22;
defparam syncload_ctrl_X22_Y16.coord_y = 16;
defparam syncload_ctrl_X22_Y16.coord_z = 1;
defparam syncload_ctrl_X22_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X22_Y19(
	.Din(),
	.Dout(SyncLoad_X22_Y19_VCC));
defparam syncload_ctrl_X22_Y19.coord_x = 19;
defparam syncload_ctrl_X22_Y19.coord_y = 17;
defparam syncload_ctrl_X22_Y19.coord_z = 1;
defparam syncload_ctrl_X22_Y19.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X22_Y8(
	.Din(),
	.Dout(SyncLoad_X22_Y8_VCC));
defparam syncload_ctrl_X22_Y8.coord_x = 10;
defparam syncload_ctrl_X22_Y8.coord_y = 17;
defparam syncload_ctrl_X22_Y8.coord_z = 1;
defparam syncload_ctrl_X22_Y8.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X23_Y15(
	.Din(),
	.Dout(SyncLoad_X23_Y15_GND));
defparam syncload_ctrl_X23_Y15.coord_x = 22;
defparam syncload_ctrl_X23_Y15.coord_y = 18;
defparam syncload_ctrl_X23_Y15.coord_z = 1;
defparam syncload_ctrl_X23_Y15.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X23_Y16(
	.Din(),
	.Dout(SyncLoad_X23_Y16_VCC));
defparam syncload_ctrl_X23_Y16.coord_x = 21;
defparam syncload_ctrl_X23_Y16.coord_y = 13;
defparam syncload_ctrl_X23_Y16.coord_z = 1;
defparam syncload_ctrl_X23_Y16.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X23_Y18(
	.Din(),
	.Dout(SyncLoad_X23_Y18_VCC));
defparam syncload_ctrl_X23_Y18.coord_x = 21;
defparam syncload_ctrl_X23_Y18.coord_y = 16;
defparam syncload_ctrl_X23_Y18.coord_z = 1;
defparam syncload_ctrl_X23_Y18.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X23_Y19(
	.Din(),
	.Dout(SyncLoad_X23_Y19_VCC));
defparam syncload_ctrl_X23_Y19.coord_x = 21;
defparam syncload_ctrl_X23_Y19.coord_y = 17;
defparam syncload_ctrl_X23_Y19.coord_z = 1;
defparam syncload_ctrl_X23_Y19.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X23_Y8(
	.Din(),
	.Dout(SyncLoad_X23_Y8_GND));
defparam syncload_ctrl_X23_Y8.coord_x = 11;
defparam syncload_ctrl_X23_Y8.coord_y = 17;
defparam syncload_ctrl_X23_Y8.coord_z = 1;
defparam syncload_ctrl_X23_Y8.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X24_Y16(
	.Din(),
	.Dout(SyncLoad_X24_Y16_GND));
defparam syncload_ctrl_X24_Y16.coord_x = 22;
defparam syncload_ctrl_X24_Y16.coord_y = 14;
defparam syncload_ctrl_X24_Y16.coord_z = 1;
defparam syncload_ctrl_X24_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X28_Y14(
	.Din(\eth_udp_inst|ip_send_inst|Equal1~1_combout ),
	.Dout(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y14_SIG ));
defparam syncload_ctrl_X28_Y14.coord_x = 21;
defparam syncload_ctrl_X28_Y14.coord_y = 9;
defparam syncload_ctrl_X28_Y14.coord_z = 1;
defparam syncload_ctrl_X28_Y14.SyncCtrlMux = 2'b10;

alta_syncctrl syncload_ctrl_X28_Y15(
	.Din(\eth_udp_inst|ip_send_inst|Equal1~1_combout ),
	.Dout(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X28_Y15_SIG ));
defparam syncload_ctrl_X28_Y15.coord_x = 21;
defparam syncload_ctrl_X28_Y15.coord_y = 10;
defparam syncload_ctrl_X28_Y15.coord_z = 1;
defparam syncload_ctrl_X28_Y15.SyncCtrlMux = 2'b10;

alta_syncctrl syncload_ctrl_X2_Y7(
	.Din(),
	.Dout(SyncLoad_X2_Y7_GND));
defparam syncload_ctrl_X2_Y7.coord_x = 9;
defparam syncload_ctrl_X2_Y7.coord_y = 12;
defparam syncload_ctrl_X2_Y7.coord_z = 1;
defparam syncload_ctrl_X2_Y7.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X4_Y7(
	.Din(),
	.Dout(SyncLoad_X4_Y7_VCC));
defparam syncload_ctrl_X4_Y7.coord_x = 17;
defparam syncload_ctrl_X4_Y7.coord_y = 12;
defparam syncload_ctrl_X4_Y7.coord_z = 1;
defparam syncload_ctrl_X4_Y7.SyncCtrlMux = 2'b01;

alta_syncctrl syncreset_ctrl_X12_Y13(
	.Din(),
	.Dout(SyncReset_X12_Y13_GND));
defparam syncreset_ctrl_X12_Y13.coord_x = 16;
defparam syncreset_ctrl_X12_Y13.coord_y = 13;
defparam syncreset_ctrl_X12_Y13.coord_z = 0;
defparam syncreset_ctrl_X12_Y13.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X12_Y14(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ));
defparam syncreset_ctrl_X12_Y14.coord_x = 2;
defparam syncreset_ctrl_X12_Y14.coord_y = 9;
defparam syncreset_ctrl_X12_Y14.coord_z = 0;
defparam syncreset_ctrl_X12_Y14.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X12_Y15(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ));
defparam syncreset_ctrl_X12_Y15.coord_x = 2;
defparam syncreset_ctrl_X12_Y15.coord_y = 10;
defparam syncreset_ctrl_X12_Y15.coord_z = 0;
defparam syncreset_ctrl_X12_Y15.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X13_Y12(
	.Din(),
	.Dout(SyncReset_X13_Y12_GND));
defparam syncreset_ctrl_X13_Y12.coord_x = 15;
defparam syncreset_ctrl_X13_Y12.coord_y = 16;
defparam syncreset_ctrl_X13_Y12.coord_z = 0;
defparam syncreset_ctrl_X13_Y12.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X14_Y12(
	.Din(),
	.Dout(SyncReset_X14_Y12_GND));
defparam syncreset_ctrl_X14_Y12.coord_x = 17;
defparam syncreset_ctrl_X14_Y12.coord_y = 16;
defparam syncreset_ctrl_X14_Y12.coord_z = 0;
defparam syncreset_ctrl_X14_Y12.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X14_Y13(
	.Din(),
	.Dout(SyncReset_X14_Y13_GND));
defparam syncreset_ctrl_X14_Y13.coord_x = 17;
defparam syncreset_ctrl_X14_Y13.coord_y = 13;
defparam syncreset_ctrl_X14_Y13.coord_z = 0;
defparam syncreset_ctrl_X14_Y13.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X14_Y17(
	.Din(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout ),
	.Dout(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X14_Y17_INV ));
defparam syncreset_ctrl_X14_Y17.coord_x = 10;
defparam syncreset_ctrl_X14_Y17.coord_y = 15;
defparam syncreset_ctrl_X14_Y17.coord_z = 0;
defparam syncreset_ctrl_X14_Y17.SyncCtrlMux = 2'b11;

alta_syncctrl syncreset_ctrl_X16_Y11(
	.Din(),
	.Dout(SyncReset_X16_Y11_GND));
defparam syncreset_ctrl_X16_Y11.coord_x = 17;
defparam syncreset_ctrl_X16_Y11.coord_y = 15;
defparam syncreset_ctrl_X16_Y11.coord_z = 0;
defparam syncreset_ctrl_X16_Y11.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X16_Y12(
	.Din(),
	.Dout(SyncReset_X16_Y12_GND));
defparam syncreset_ctrl_X16_Y12.coord_x = 16;
defparam syncreset_ctrl_X16_Y12.coord_y = 16;
defparam syncreset_ctrl_X16_Y12.coord_z = 0;
defparam syncreset_ctrl_X16_Y12.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X16_Y13(
	.Din(),
	.Dout(SyncReset_X16_Y13_GND));
defparam syncreset_ctrl_X16_Y13.coord_x = 17;
defparam syncreset_ctrl_X16_Y13.coord_y = 14;
defparam syncreset_ctrl_X16_Y13.coord_z = 0;
defparam syncreset_ctrl_X16_Y13.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X17_Y13(
	.Din(),
	.Dout(SyncReset_X17_Y13_GND));
defparam syncreset_ctrl_X17_Y13.coord_x = 16;
defparam syncreset_ctrl_X17_Y13.coord_y = 15;
defparam syncreset_ctrl_X17_Y13.coord_z = 0;
defparam syncreset_ctrl_X17_Y13.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X1_Y17(
	.Din(\camera_if_inst|cam_vsync_r [0]),
	.Dout(\camera_if_inst|cam_vsync_r[0]__SyncReset_X1_Y17_SIG ));
defparam syncreset_ctrl_X1_Y17.coord_x = 11;
defparam syncreset_ctrl_X1_Y17.coord_y = 16;
defparam syncreset_ctrl_X1_Y17.coord_z = 0;
defparam syncreset_ctrl_X1_Y17.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X1_Y7(
	.Din(),
	.Dout(SyncReset_X1_Y7_GND));
defparam syncreset_ctrl_X1_Y7.coord_x = 8;
defparam syncreset_ctrl_X1_Y7.coord_y = 12;
defparam syncreset_ctrl_X1_Y7.coord_z = 0;
defparam syncreset_ctrl_X1_Y7.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X22_Y16(
	.Din(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Dout(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X22_Y16_SIG ));
defparam syncreset_ctrl_X22_Y16.coord_x = 22;
defparam syncreset_ctrl_X22_Y16.coord_y = 16;
defparam syncreset_ctrl_X22_Y16.coord_z = 0;
defparam syncreset_ctrl_X22_Y16.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X22_Y19(
	.Din(),
	.Dout(SyncReset_X22_Y19_GND));
defparam syncreset_ctrl_X22_Y19.coord_x = 19;
defparam syncreset_ctrl_X22_Y19.coord_y = 17;
defparam syncreset_ctrl_X22_Y19.coord_z = 0;
defparam syncreset_ctrl_X22_Y19.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X22_Y8(
	.Din(),
	.Dout(SyncReset_X22_Y8_GND));
defparam syncreset_ctrl_X22_Y8.coord_x = 10;
defparam syncreset_ctrl_X22_Y8.coord_y = 17;
defparam syncreset_ctrl_X22_Y8.coord_z = 0;
defparam syncreset_ctrl_X22_Y8.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X23_Y15(
	.Din(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Dout(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X23_Y15_SIG ));
defparam syncreset_ctrl_X23_Y15.coord_x = 22;
defparam syncreset_ctrl_X23_Y15.coord_y = 18;
defparam syncreset_ctrl_X23_Y15.coord_z = 0;
defparam syncreset_ctrl_X23_Y15.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X23_Y16(
	.Din(),
	.Dout(SyncReset_X23_Y16_GND));
defparam syncreset_ctrl_X23_Y16.coord_x = 21;
defparam syncreset_ctrl_X23_Y16.coord_y = 13;
defparam syncreset_ctrl_X23_Y16.coord_z = 0;
defparam syncreset_ctrl_X23_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X23_Y18(
	.Din(),
	.Dout(SyncReset_X23_Y18_GND));
defparam syncreset_ctrl_X23_Y18.coord_x = 21;
defparam syncreset_ctrl_X23_Y18.coord_y = 16;
defparam syncreset_ctrl_X23_Y18.coord_z = 0;
defparam syncreset_ctrl_X23_Y18.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X23_Y19(
	.Din(),
	.Dout(SyncReset_X23_Y19_GND));
defparam syncreset_ctrl_X23_Y19.coord_x = 21;
defparam syncreset_ctrl_X23_Y19.coord_y = 17;
defparam syncreset_ctrl_X23_Y19.coord_z = 0;
defparam syncreset_ctrl_X23_Y19.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X23_Y8(
	.Din(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout ),
	.Dout(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X23_Y8_INV ));
defparam syncreset_ctrl_X23_Y8.coord_x = 11;
defparam syncreset_ctrl_X23_Y8.coord_y = 17;
defparam syncreset_ctrl_X23_Y8.coord_z = 0;
defparam syncreset_ctrl_X23_Y8.SyncCtrlMux = 2'b11;

alta_syncctrl syncreset_ctrl_X24_Y16(
	.Din(\eth_udp_inst|ip_send_inst|cnt[3]~11_combout ),
	.Dout(\eth_udp_inst|ip_send_inst|cnt[3]~11_combout__SyncReset_X24_Y16_SIG ));
defparam syncreset_ctrl_X24_Y16.coord_x = 22;
defparam syncreset_ctrl_X24_Y16.coord_y = 14;
defparam syncreset_ctrl_X24_Y16.coord_z = 0;
defparam syncreset_ctrl_X24_Y16.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X28_Y14(
	.Din(),
	.Dout(SyncReset_X28_Y14_GND));
defparam syncreset_ctrl_X28_Y14.coord_x = 21;
defparam syncreset_ctrl_X28_Y14.coord_y = 9;
defparam syncreset_ctrl_X28_Y14.coord_z = 0;
defparam syncreset_ctrl_X28_Y14.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X28_Y15(
	.Din(),
	.Dout(SyncReset_X28_Y15_GND));
defparam syncreset_ctrl_X28_Y15.coord_x = 21;
defparam syncreset_ctrl_X28_Y15.coord_y = 10;
defparam syncreset_ctrl_X28_Y15.coord_z = 0;
defparam syncreset_ctrl_X28_Y15.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X2_Y7(
	.Din(\camera_if_inst|cam_hsync_r [0]),
	.Dout(\camera_if_inst|cam_hsync_r[0]__SyncReset_X2_Y7_INV ));
defparam syncreset_ctrl_X2_Y7.coord_x = 9;
defparam syncreset_ctrl_X2_Y7.coord_y = 12;
defparam syncreset_ctrl_X2_Y7.coord_z = 0;
defparam syncreset_ctrl_X2_Y7.SyncCtrlMux = 2'b11;

alta_syncctrl syncreset_ctrl_X4_Y7(
	.Din(),
	.Dout(SyncReset_X4_Y7_GND));
defparam syncreset_ctrl_X4_Y7.coord_x = 17;
defparam syncreset_ctrl_X4_Y7.coord_y = 12;
defparam syncreset_ctrl_X4_Y7.coord_z = 0;
defparam syncreset_ctrl_X4_Y7.SyncCtrlMux = 2'b00;

alta_slice \timer[0] (
	.A(vcc),
	.B(timer[0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(timer[0]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y15_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y15_GND),
	.LutOut(\timer[0]~25_combout ),
	.Cout(\timer[0]~26 ),
	.Q(timer[0]));
defparam \timer[0] .coord_x = 2;
defparam \timer[0] .coord_y = 10;
defparam \timer[0] .coord_z = 4;
defparam \timer[0] .mask = 16'h33CC;
defparam \timer[0] .modeMux = 1'b0;
defparam \timer[0] .FeedbackMux = 1'b0;
defparam \timer[0] .ShiftMux = 1'b0;
defparam \timer[0] .BypassEn = 1'b1;
defparam \timer[0] .CarryEnb = 1'b0;

alta_slice \timer[10] (
	.A(vcc),
	.B(timer[10]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[9]~44 ),
	.Qin(timer[10]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y15_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y15_GND),
	.LutOut(\timer[10]~45_combout ),
	.Cout(\timer[10]~46 ),
	.Q(timer[10]));
defparam \timer[10] .coord_x = 2;
defparam \timer[10] .coord_y = 10;
defparam \timer[10] .coord_z = 14;
defparam \timer[10] .mask = 16'hC30C;
defparam \timer[10] .modeMux = 1'b1;
defparam \timer[10] .FeedbackMux = 1'b0;
defparam \timer[10] .ShiftMux = 1'b0;
defparam \timer[10] .BypassEn = 1'b1;
defparam \timer[10] .CarryEnb = 1'b0;

alta_slice \timer[11] (
	.A(timer[11]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[10]~46 ),
	.Qin(timer[11]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y15_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y15_GND),
	.LutOut(\timer[11]~47_combout ),
	.Cout(\timer[11]~48 ),
	.Q(timer[11]));
defparam \timer[11] .coord_x = 2;
defparam \timer[11] .coord_y = 10;
defparam \timer[11] .coord_z = 15;
defparam \timer[11] .mask = 16'h5A5F;
defparam \timer[11] .modeMux = 1'b1;
defparam \timer[11] .FeedbackMux = 1'b0;
defparam \timer[11] .ShiftMux = 1'b0;
defparam \timer[11] .BypassEn = 1'b1;
defparam \timer[11] .CarryEnb = 1'b0;

alta_slice \timer[12] (
	.A(vcc),
	.B(timer[12]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[11]~48 ),
	.Qin(timer[12]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_GND),
	.LutOut(\timer[12]~49_combout ),
	.Cout(\timer[12]~50 ),
	.Q(timer[12]));
defparam \timer[12] .coord_x = 2;
defparam \timer[12] .coord_y = 9;
defparam \timer[12] .coord_z = 0;
defparam \timer[12] .mask = 16'hC30C;
defparam \timer[12] .modeMux = 1'b1;
defparam \timer[12] .FeedbackMux = 1'b0;
defparam \timer[12] .ShiftMux = 1'b0;
defparam \timer[12] .BypassEn = 1'b1;
defparam \timer[12] .CarryEnb = 1'b0;

alta_slice \timer[13] (
	.A(timer[13]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[12]~50 ),
	.Qin(timer[13]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_GND),
	.LutOut(\timer[13]~51_combout ),
	.Cout(\timer[13]~52 ),
	.Q(timer[13]));
defparam \timer[13] .coord_x = 2;
defparam \timer[13] .coord_y = 9;
defparam \timer[13] .coord_z = 1;
defparam \timer[13] .mask = 16'h5A5F;
defparam \timer[13] .modeMux = 1'b1;
defparam \timer[13] .FeedbackMux = 1'b0;
defparam \timer[13] .ShiftMux = 1'b0;
defparam \timer[13] .BypassEn = 1'b1;
defparam \timer[13] .CarryEnb = 1'b0;

alta_slice \timer[14] (
	.A(vcc),
	.B(timer[14]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[13]~52 ),
	.Qin(timer[14]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_GND),
	.LutOut(\timer[14]~53_combout ),
	.Cout(\timer[14]~54 ),
	.Q(timer[14]));
defparam \timer[14] .coord_x = 2;
defparam \timer[14] .coord_y = 9;
defparam \timer[14] .coord_z = 2;
defparam \timer[14] .mask = 16'hC30C;
defparam \timer[14] .modeMux = 1'b1;
defparam \timer[14] .FeedbackMux = 1'b0;
defparam \timer[14] .ShiftMux = 1'b0;
defparam \timer[14] .BypassEn = 1'b1;
defparam \timer[14] .CarryEnb = 1'b0;

alta_slice \timer[15] (
	.A(timer[15]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[14]~54 ),
	.Qin(timer[15]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_GND),
	.LutOut(\timer[15]~55_combout ),
	.Cout(\timer[15]~56 ),
	.Q(timer[15]));
defparam \timer[15] .coord_x = 2;
defparam \timer[15] .coord_y = 9;
defparam \timer[15] .coord_z = 3;
defparam \timer[15] .mask = 16'h5A5F;
defparam \timer[15] .modeMux = 1'b1;
defparam \timer[15] .FeedbackMux = 1'b0;
defparam \timer[15] .ShiftMux = 1'b0;
defparam \timer[15] .BypassEn = 1'b1;
defparam \timer[15] .CarryEnb = 1'b0;

alta_slice \timer[16] (
	.A(timer[16]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[15]~56 ),
	.Qin(timer[16]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_GND),
	.LutOut(\timer[16]~57_combout ),
	.Cout(\timer[16]~58 ),
	.Q(timer[16]));
defparam \timer[16] .coord_x = 2;
defparam \timer[16] .coord_y = 9;
defparam \timer[16] .coord_z = 4;
defparam \timer[16] .mask = 16'hA50A;
defparam \timer[16] .modeMux = 1'b1;
defparam \timer[16] .FeedbackMux = 1'b0;
defparam \timer[16] .ShiftMux = 1'b0;
defparam \timer[16] .BypassEn = 1'b1;
defparam \timer[16] .CarryEnb = 1'b0;

alta_slice \timer[17] (
	.A(timer[17]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[16]~58 ),
	.Qin(timer[17]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_GND),
	.LutOut(\timer[17]~59_combout ),
	.Cout(\timer[17]~60 ),
	.Q(timer[17]));
defparam \timer[17] .coord_x = 2;
defparam \timer[17] .coord_y = 9;
defparam \timer[17] .coord_z = 5;
defparam \timer[17] .mask = 16'h5A5F;
defparam \timer[17] .modeMux = 1'b1;
defparam \timer[17] .FeedbackMux = 1'b0;
defparam \timer[17] .ShiftMux = 1'b0;
defparam \timer[17] .BypassEn = 1'b1;
defparam \timer[17] .CarryEnb = 1'b0;

alta_slice \timer[18] (
	.A(vcc),
	.B(timer[18]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[17]~60 ),
	.Qin(timer[18]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_GND),
	.LutOut(\timer[18]~61_combout ),
	.Cout(\timer[18]~62 ),
	.Q(timer[18]));
defparam \timer[18] .coord_x = 2;
defparam \timer[18] .coord_y = 9;
defparam \timer[18] .coord_z = 6;
defparam \timer[18] .mask = 16'hC30C;
defparam \timer[18] .modeMux = 1'b1;
defparam \timer[18] .FeedbackMux = 1'b0;
defparam \timer[18] .ShiftMux = 1'b0;
defparam \timer[18] .BypassEn = 1'b1;
defparam \timer[18] .CarryEnb = 1'b0;

alta_slice \timer[19] (
	.A(vcc),
	.B(timer[19]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[18]~62 ),
	.Qin(timer[19]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_GND),
	.LutOut(\timer[19]~63_combout ),
	.Cout(\timer[19]~64 ),
	.Q(timer[19]));
defparam \timer[19] .coord_x = 2;
defparam \timer[19] .coord_y = 9;
defparam \timer[19] .coord_z = 7;
defparam \timer[19] .mask = 16'h3C3F;
defparam \timer[19] .modeMux = 1'b1;
defparam \timer[19] .FeedbackMux = 1'b0;
defparam \timer[19] .ShiftMux = 1'b0;
defparam \timer[19] .BypassEn = 1'b1;
defparam \timer[19] .CarryEnb = 1'b0;

alta_slice \timer[1] (
	.A(timer[1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[0]~26 ),
	.Qin(timer[1]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y15_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y15_GND),
	.LutOut(\timer[1]~27_combout ),
	.Cout(\timer[1]~28 ),
	.Q(timer[1]));
defparam \timer[1] .coord_x = 2;
defparam \timer[1] .coord_y = 10;
defparam \timer[1] .coord_z = 5;
defparam \timer[1] .mask = 16'h5A5F;
defparam \timer[1] .modeMux = 1'b1;
defparam \timer[1] .FeedbackMux = 1'b0;
defparam \timer[1] .ShiftMux = 1'b0;
defparam \timer[1] .BypassEn = 1'b1;
defparam \timer[1] .CarryEnb = 1'b0;

alta_slice \timer[20] (
	.A(vcc),
	.B(timer[20]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[19]~64 ),
	.Qin(timer[20]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_GND),
	.LutOut(\timer[20]~65_combout ),
	.Cout(\timer[20]~66 ),
	.Q(timer[20]));
defparam \timer[20] .coord_x = 2;
defparam \timer[20] .coord_y = 9;
defparam \timer[20] .coord_z = 8;
defparam \timer[20] .mask = 16'hC30C;
defparam \timer[20] .modeMux = 1'b1;
defparam \timer[20] .FeedbackMux = 1'b0;
defparam \timer[20] .ShiftMux = 1'b0;
defparam \timer[20] .BypassEn = 1'b1;
defparam \timer[20] .CarryEnb = 1'b0;

alta_slice \timer[21] (
	.A(timer[21]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[20]~66 ),
	.Qin(timer[21]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_GND),
	.LutOut(\timer[21]~67_combout ),
	.Cout(\timer[21]~68 ),
	.Q(timer[21]));
defparam \timer[21] .coord_x = 2;
defparam \timer[21] .coord_y = 9;
defparam \timer[21] .coord_z = 9;
defparam \timer[21] .mask = 16'h5A5F;
defparam \timer[21] .modeMux = 1'b1;
defparam \timer[21] .FeedbackMux = 1'b0;
defparam \timer[21] .ShiftMux = 1'b0;
defparam \timer[21] .BypassEn = 1'b1;
defparam \timer[21] .CarryEnb = 1'b0;

alta_slice \timer[22] (
	.A(vcc),
	.B(timer[22]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[21]~68 ),
	.Qin(timer[22]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_GND),
	.LutOut(\timer[22]~69_combout ),
	.Cout(\timer[22]~70 ),
	.Q(timer[22]));
defparam \timer[22] .coord_x = 2;
defparam \timer[22] .coord_y = 9;
defparam \timer[22] .coord_z = 10;
defparam \timer[22] .mask = 16'hC30C;
defparam \timer[22] .modeMux = 1'b1;
defparam \timer[22] .FeedbackMux = 1'b0;
defparam \timer[22] .ShiftMux = 1'b0;
defparam \timer[22] .BypassEn = 1'b1;
defparam \timer[22] .CarryEnb = 1'b0;

alta_slice \timer[23] (
	.A(timer[23]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[22]~70 ),
	.Qin(timer[23]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_GND),
	.LutOut(\timer[23]~71_combout ),
	.Cout(\timer[23]~72 ),
	.Q(timer[23]));
defparam \timer[23] .coord_x = 2;
defparam \timer[23] .coord_y = 9;
defparam \timer[23] .coord_z = 11;
defparam \timer[23] .mask = 16'h5A5F;
defparam \timer[23] .modeMux = 1'b1;
defparam \timer[23] .FeedbackMux = 1'b0;
defparam \timer[23] .ShiftMux = 1'b0;
defparam \timer[23] .BypassEn = 1'b1;
defparam \timer[23] .CarryEnb = 1'b0;

alta_slice \timer[24] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(timer[24]),
	.Cin(\timer[23]~72 ),
	.Qin(timer[24]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y14_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_GND),
	.LutOut(\timer[24]~73_combout ),
	.Cout(),
	.Q(timer[24]));
defparam \timer[24] .coord_x = 2;
defparam \timer[24] .coord_y = 9;
defparam \timer[24] .coord_z = 12;
defparam \timer[24] .mask = 16'hF00F;
defparam \timer[24] .modeMux = 1'b1;
defparam \timer[24] .FeedbackMux = 1'b0;
defparam \timer[24] .ShiftMux = 1'b0;
defparam \timer[24] .BypassEn = 1'b1;
defparam \timer[24] .CarryEnb = 1'b1;

alta_slice \timer[2] (
	.A(timer[2]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[1]~28 ),
	.Qin(timer[2]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y15_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y15_GND),
	.LutOut(\timer[2]~29_combout ),
	.Cout(\timer[2]~30 ),
	.Q(timer[2]));
defparam \timer[2] .coord_x = 2;
defparam \timer[2] .coord_y = 10;
defparam \timer[2] .coord_z = 6;
defparam \timer[2] .mask = 16'hA50A;
defparam \timer[2] .modeMux = 1'b1;
defparam \timer[2] .FeedbackMux = 1'b0;
defparam \timer[2] .ShiftMux = 1'b0;
defparam \timer[2] .BypassEn = 1'b1;
defparam \timer[2] .CarryEnb = 1'b0;

alta_slice \timer[3] (
	.A(vcc),
	.B(timer[3]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[2]~30 ),
	.Qin(timer[3]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y15_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y15_GND),
	.LutOut(\timer[3]~31_combout ),
	.Cout(\timer[3]~32 ),
	.Q(timer[3]));
defparam \timer[3] .coord_x = 2;
defparam \timer[3] .coord_y = 10;
defparam \timer[3] .coord_z = 7;
defparam \timer[3] .mask = 16'h3C3F;
defparam \timer[3] .modeMux = 1'b1;
defparam \timer[3] .FeedbackMux = 1'b0;
defparam \timer[3] .ShiftMux = 1'b0;
defparam \timer[3] .BypassEn = 1'b1;
defparam \timer[3] .CarryEnb = 1'b0;

alta_slice \timer[4] (
	.A(vcc),
	.B(timer[4]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[3]~32 ),
	.Qin(timer[4]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y15_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y15_GND),
	.LutOut(\timer[4]~33_combout ),
	.Cout(\timer[4]~34 ),
	.Q(timer[4]));
defparam \timer[4] .coord_x = 2;
defparam \timer[4] .coord_y = 10;
defparam \timer[4] .coord_z = 8;
defparam \timer[4] .mask = 16'hC30C;
defparam \timer[4] .modeMux = 1'b1;
defparam \timer[4] .FeedbackMux = 1'b0;
defparam \timer[4] .ShiftMux = 1'b0;
defparam \timer[4] .BypassEn = 1'b1;
defparam \timer[4] .CarryEnb = 1'b0;

alta_slice \timer[5] (
	.A(vcc),
	.B(timer[5]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[4]~34 ),
	.Qin(timer[5]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y15_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y15_GND),
	.LutOut(\timer[5]~35_combout ),
	.Cout(\timer[5]~36 ),
	.Q(timer[5]));
defparam \timer[5] .coord_x = 2;
defparam \timer[5] .coord_y = 10;
defparam \timer[5] .coord_z = 9;
defparam \timer[5] .mask = 16'h3C3F;
defparam \timer[5] .modeMux = 1'b1;
defparam \timer[5] .FeedbackMux = 1'b0;
defparam \timer[5] .ShiftMux = 1'b0;
defparam \timer[5] .BypassEn = 1'b1;
defparam \timer[5] .CarryEnb = 1'b0;

alta_slice \timer[6] (
	.A(vcc),
	.B(timer[6]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[5]~36 ),
	.Qin(timer[6]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y15_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y15_GND),
	.LutOut(\timer[6]~37_combout ),
	.Cout(\timer[6]~38 ),
	.Q(timer[6]));
defparam \timer[6] .coord_x = 2;
defparam \timer[6] .coord_y = 10;
defparam \timer[6] .coord_z = 10;
defparam \timer[6] .mask = 16'hC30C;
defparam \timer[6] .modeMux = 1'b1;
defparam \timer[6] .FeedbackMux = 1'b0;
defparam \timer[6] .ShiftMux = 1'b0;
defparam \timer[6] .BypassEn = 1'b1;
defparam \timer[6] .CarryEnb = 1'b0;

alta_slice \timer[7] (
	.A(timer[7]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[6]~38 ),
	.Qin(timer[7]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y15_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y15_GND),
	.LutOut(\timer[7]~39_combout ),
	.Cout(\timer[7]~40 ),
	.Q(timer[7]));
defparam \timer[7] .coord_x = 2;
defparam \timer[7] .coord_y = 10;
defparam \timer[7] .coord_z = 11;
defparam \timer[7] .mask = 16'h5A5F;
defparam \timer[7] .modeMux = 1'b1;
defparam \timer[7] .FeedbackMux = 1'b0;
defparam \timer[7] .ShiftMux = 1'b0;
defparam \timer[7] .BypassEn = 1'b1;
defparam \timer[7] .CarryEnb = 1'b0;

alta_slice \timer[8] (
	.A(timer[8]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[7]~40 ),
	.Qin(timer[8]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y15_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y15_GND),
	.LutOut(\timer[8]~41_combout ),
	.Cout(\timer[8]~42 ),
	.Q(timer[8]));
defparam \timer[8] .coord_x = 2;
defparam \timer[8] .coord_y = 10;
defparam \timer[8] .coord_z = 12;
defparam \timer[8] .mask = 16'hA50A;
defparam \timer[8] .modeMux = 1'b1;
defparam \timer[8] .FeedbackMux = 1'b0;
defparam \timer[8] .ShiftMux = 1'b0;
defparam \timer[8] .BypassEn = 1'b1;
defparam \timer[8] .CarryEnb = 1'b0;

alta_slice \timer[9] (
	.A(vcc),
	.B(timer[9]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[8]~42 ),
	.Qin(timer[9]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y15_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X12_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y15_GND),
	.LutOut(\timer[9]~43_combout ),
	.Cout(\timer[9]~44 ),
	.Q(timer[9]));
defparam \timer[9] .coord_x = 2;
defparam \timer[9] .coord_y = 10;
defparam \timer[9] .coord_z = 13;
defparam \timer[9] .mask = 16'h3C3F;
defparam \timer[9] .modeMux = 1'b1;
defparam \timer[9] .FeedbackMux = 1'b0;
defparam \timer[9] .ShiftMux = 1'b0;
defparam \timer[9] .BypassEn = 1'b1;
defparam \timer[9] .CarryEnb = 1'b0;

endmodule
