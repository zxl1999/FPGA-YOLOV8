`timescale 1 ps/ 1 ps

module top_fpga(
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	clk,
	rst_n,
	cam_scl,
	cam_sda,
	cam_data,
	cam_vsync,
	cam_hsync,
	cam_pclk,
	cam_xclk,
	cam_pdown,
	cam_reset,
	e_txen,
	e_tx,
	e_rxer,
	e_rxdv,
	e_rxclk,
	e_rx,
	led);
input	altera_reserved_tms;
input	altera_reserved_tck;
input	altera_reserved_tdi;
output	altera_reserved_tdo;
input	clk;
input	rst_n;
output	cam_scl;
inout	cam_sda;
input	[7:0] cam_data;
input	cam_vsync;
input	cam_hsync;
input	cam_pclk;
output	cam_xclk;
output	cam_pdown;
output	cam_reset;
output	e_txen;
output	[1:0] e_tx;
input	e_rxer;
input	e_rxdv;
input	e_rxclk;
input	[1:0] e_rx;
output	led;

//wire	gnd;
//wire	vcc;
wire	\Add0~0_combout ;
wire	\Add0~1 ;
wire	\Add0~2_combout ;
wire	\Add0~3 ;
wire	\Add0~4_combout ;
wire	\Add0~5 ;
wire	\Add0~6_combout ;
wire	\Add0~7 ;
wire	\Add0~8_combout ;
wire	AsyncReset_X11_Y14_GND;
wire	AsyncReset_X11_Y16_GND;
wire	AsyncReset_X12_Y14_GND;
wire	AsyncReset_X12_Y16_GND;
wire	AsyncReset_X12_Y18_GND;
wire	AsyncReset_X13_Y16_GND;
wire	AsyncReset_X13_Y18_GND;
wire	AsyncReset_X14_Y14_GND;
wire	AsyncReset_X14_Y16_GND;
wire	AsyncReset_X14_Y18_GND;
wire	AsyncReset_X14_Y19_GND;
wire	AsyncReset_X14_Y20_GND;
wire	AsyncReset_X16_Y10_GND;
wire	AsyncReset_X16_Y12_GND;
wire	AsyncReset_X16_Y16_GND;
wire	AsyncReset_X16_Y17_GND;
wire	AsyncReset_X16_Y18_GND;
wire	AsyncReset_X16_Y19_GND;
wire	AsyncReset_X16_Y8_GND;
wire	AsyncReset_X17_Y15_GND;
wire	AsyncReset_X17_Y16_GND;
wire	AsyncReset_X17_Y18_GND;
wire	AsyncReset_X17_Y19_GND;
wire	AsyncReset_X17_Y20_GND;
wire	AsyncReset_X18_Y13_GND;
wire	AsyncReset_X18_Y15_GND;
wire	AsyncReset_X18_Y16_GND;
wire	AsyncReset_X18_Y18_GND;
wire	AsyncReset_X18_Y19_GND;
wire	AsyncReset_X18_Y20_GND;
wire	AsyncReset_X19_Y16_GND;
wire	AsyncReset_X19_Y18_GND;
wire	AsyncReset_X19_Y19_GND;
wire	AsyncReset_X1_Y7_GND;
wire	AsyncReset_X21_Y15_GND;
wire	AsyncReset_X21_Y17_GND;
wire	AsyncReset_X21_Y18_GND;
wire	AsyncReset_X21_Y20_GND;
wire	AsyncReset_X22_Y14_GND;
wire	AsyncReset_X22_Y15_GND;
wire	AsyncReset_X22_Y17_GND;
wire	AsyncReset_X22_Y18_GND;
wire	AsyncReset_X24_Y18_GND;
wire	AsyncReset_X25_Y15_GND;
wire	AsyncReset_X25_Y18_GND;
wire	AsyncReset_X25_Y19_GND;
wire	AsyncReset_X2_Y7_GND;
wire	AsyncReset_X33_Y12_GND;
wire	AsyncReset_X5_Y7_GND;
wire	AsyncReset_X9_Y7_GND;
wire	\Equal0~0_combout ;
wire	\Equal0~1_combout ;
wire	\Equal0~2_combout ;
wire	\Equal0~3_combout ;
wire	\Equal0~4_combout ;
wire	\Equal0~5_combout ;
wire	\Equal0~6_combout ;
wire	\Equal0~7_combout ;
wire	\LessThan0~0_combout ;
wire	SyncLoad_X10_Y9_VCC;
wire	SyncLoad_X11_Y14_VCC;
wire	SyncLoad_X11_Y16_VCC;
wire	SyncLoad_X11_Y9_VCC;
wire	SyncLoad_X12_Y14_VCC;
wire	SyncLoad_X12_Y16_VCC;
wire	SyncLoad_X12_Y18_VCC;
wire	SyncLoad_X13_Y10_VCC;
wire	SyncLoad_X13_Y16_VCC;
wire	SyncLoad_X13_Y18_VCC;
wire	SyncLoad_X13_Y7_VCC;
wire	SyncLoad_X14_Y10_VCC;
wire	SyncLoad_X14_Y16_VCC;
wire	SyncLoad_X14_Y18_VCC;
wire	SyncLoad_X14_Y8_VCC;
wire	SyncLoad_X14_Y9_VCC;
wire	SyncLoad_X16_Y14_VCC;
wire	SyncLoad_X16_Y16_VCC;
wire	SyncLoad_X16_Y18_VCC;
wire	SyncLoad_X16_Y19_VCC;
wire	SyncLoad_X16_Y9_VCC;
wire	SyncLoad_X17_Y15_GND;
wire	SyncLoad_X17_Y17_VCC;
wire	SyncLoad_X17_Y9_VCC;
wire	SyncLoad_X18_Y13_GND;
wire	SyncLoad_X18_Y15_GND;
wire	SyncLoad_X18_Y17_VCC;
wire	SyncLoad_X18_Y19_VCC;
wire	SyncLoad_X19_Y16_VCC;
wire	SyncLoad_X19_Y17_VCC;
wire	SyncLoad_X19_Y8_GND;
wire	SyncLoad_X1_Y7_GND;
wire	SyncLoad_X21_Y15_GND;
wire	SyncLoad_X21_Y17_GND;
wire	SyncLoad_X21_Y18_VCC;
wire	SyncLoad_X21_Y19_VCC;
wire	SyncLoad_X23_Y16_VCC;
wire	SyncLoad_X24_Y15_GND;
wire	SyncLoad_X24_Y16_VCC;
wire	SyncLoad_X24_Y19_VCC;
wire	SyncLoad_X25_Y12_VCC;
wire	SyncLoad_X25_Y18_GND;
wire	SyncLoad_X25_Y19_GND;
wire	SyncLoad_X26_Y15_GND;
wire	SyncLoad_X26_Y16_GND;
wire	SyncLoad_X28_Y9_VCC;
wire	SyncLoad_X29_Y9_GND;
wire	SyncLoad_X2_Y7_VCC;
wire	SyncLoad_X33_Y16_VCC;
wire	SyncLoad_X5_Y7_GND;
wire	SyncLoad_X9_Y7_VCC;
wire	SyncReset_X10_Y9_GND;
wire	SyncReset_X11_Y14_GND;
wire	SyncReset_X11_Y16_GND;
wire	SyncReset_X11_Y9_GND;
wire	SyncReset_X12_Y14_GND;
wire	SyncReset_X12_Y16_GND;
wire	SyncReset_X12_Y18_GND;
wire	SyncReset_X13_Y10_GND;
wire	SyncReset_X13_Y16_GND;
wire	SyncReset_X13_Y18_GND;
wire	SyncReset_X13_Y7_GND;
wire	SyncReset_X14_Y10_GND;
wire	SyncReset_X14_Y16_GND;
wire	SyncReset_X14_Y18_GND;
wire	SyncReset_X14_Y8_GND;
wire	SyncReset_X14_Y9_GND;
wire	SyncReset_X16_Y14_GND;
wire	SyncReset_X16_Y16_GND;
wire	SyncReset_X16_Y17_GND;
wire	SyncReset_X16_Y18_GND;
wire	SyncReset_X16_Y19_GND;
wire	SyncReset_X16_Y9_GND;
wire	SyncReset_X17_Y16_GND;
wire	SyncReset_X17_Y17_GND;
wire	SyncReset_X17_Y20_GND;
wire	SyncReset_X17_Y9_GND;
wire	SyncReset_X18_Y16_GND;
wire	SyncReset_X18_Y17_GND;
wire	SyncReset_X18_Y18_GND;
wire	SyncReset_X18_Y19_GND;
wire	SyncReset_X18_Y20_GND;
wire	SyncReset_X19_Y16_GND;
wire	SyncReset_X19_Y17_GND;
wire	SyncReset_X21_Y16_GND;
wire	SyncReset_X21_Y18_GND;
wire	SyncReset_X21_Y19_GND;
wire	SyncReset_X22_Y14_GND;
wire	SyncReset_X22_Y15_GND;
wire	SyncReset_X23_Y16_GND;
wire	SyncReset_X24_Y16_GND;
wire	SyncReset_X24_Y19_GND;
wire	SyncReset_X25_Y12_GND;
wire	SyncReset_X28_Y9_GND;
wire	SyncReset_X2_Y7_GND;
wire	SyncReset_X33_Y16_GND;
wire	SyncReset_X9_Y7_GND;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y11_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y10_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y11_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y10_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y11_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X19_Y8_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y14_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y15_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y12_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y12_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y13_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y15_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y12_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y13_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y16_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y9_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~combout ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ;
wire	[4:0] \alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus ;
//wire	\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [0];
//wire	\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [1];
//wire	\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [2];
//wire	\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [3];
//wire	\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [4];
wire	\alt_pll_inst|altpll_component|auto_generated|pll_lock_sync~feeder_combout ;
wire	\alt_pll_inst|altpll_component|auto_generated|pll_lock_sync~q ;
wire	[4:0] \alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk ;
//wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk [0];
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X17_Y11_SIG_VCC ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X28_Y9_SIG_VCC ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X16_Y11_SIG_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y11_SIG_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y10_SIG_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y11_SIG_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y10_SIG_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y11_SIG_SIG ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X19_Y8_SIG_SIG ;
//wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk [1];
//wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk [2];
//wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk [3];
//wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk [4];
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_fbout ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked ;
wire	\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked_X1_Y1_SIG_VCC ;
wire	\altera_internal_jtag~TCKUTAP ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y14_SIG_VCC ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y15_SIG_VCC ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y17_SIG_VCC ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y18_SIG_VCC ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y19_SIG_VCC ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y20_SIG_VCC ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y13_SIG_VCC ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y18_SIG_VCC ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y15_SIG_VCC ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y17_SIG_VCC ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y18_SIG_VCC ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout_X18_Y13_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout_X18_Y16_INV_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout_X18_Y16_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17_combout_X17_Y15_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17_combout_X18_Y15_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20_combout_X18_Y15_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout_X19_Y16_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout_X19_Y16_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X17_Y17_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X18_Y17_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y18_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y19_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X18_Y20_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout_X18_Y17_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout_X17_Y16_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11]_X19_Y17_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout_X19_Y17_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q_X21_Y16_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12_combout_X22_Y17_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10_combout_X22_Y17_SIG_INV ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X18_Y18_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0_combout_X18_Y20_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena~combout_X16_Y17_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X19_Y18_SIG_INV ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X22_Y18_SIG_INV ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X19_Y18_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X22_Y18_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X11_Y14_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y14_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y18_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X13_Y18_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ;
wire	\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X24_Y19_SIG_SIG ;
wire	\altera_internal_jtag~TDIUTAP ;
wire	\altera_internal_jtag~TDO ;
wire	\altera_internal_jtag~TMSUTAP ;
wire	\altera_internal_jtag~TMSUTAP__SyncReset_X17_Y15_SIG ;
wire	\altera_internal_jtag~TMSUTAP__SyncReset_X18_Y13_SIG ;
wire	\altera_internal_jtag~TMSUTAP__SyncReset_X21_Y15_INV ;
wire	\altera_internal_jtag~TMSUTAP__SyncReset_X21_Y17_SIG ;
wire	\altera_reserved_tck~input_o ;
wire	\altera_reserved_tdi~input_o ;
wire	\altera_reserved_tms~input_o ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X17_Y15_SIG ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X17_Y17_SIG ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X21_Y16_SIG ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout__SyncLoad_X18_Y16_SIG ;
wire	[3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~16_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~24_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ;
wire	[3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~15_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~18_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ;
wire	[4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~10 ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13_combout__SyncReset_X18_Y15_SIG ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~9_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~11_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~12 ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~14_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~16_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~17 ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~18_combout ;
wire	[3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ;
wire	[2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ;
wire	[3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ;
wire	[3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5]~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~feeder_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~feeder_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8]~feeder_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8]~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9]~feeder_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9]~q ;
wire	[10:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~6_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~7_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~8_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~9_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [6];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [7];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [8];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [9];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~10_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~11_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~12_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~13_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~14_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~15_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~3_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~4_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ;
wire	[9:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9];
wire	[4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~8 ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~11_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~12 ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~14 ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~16 ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout__SyncLoad_X17_Y16_SIG ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ;
wire	[15:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3]__SyncLoad_X21_Y16_SIG ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8]__AsyncReset_X18_Y16_SIG ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ;
wire	[2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt ;
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1];
//wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2];
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ;
wire	\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q__AsyncReset_X18_Y13_INV ;
wire	\auto_hub|~GND~combout ;
wire	[7:0] \auto_signaltap_0|acq_data_in_reg ;
//wire	\auto_signaltap_0|acq_data_in_reg [0];
wire	\auto_signaltap_0|acq_data_in_reg[0]~feeder_combout ;
//wire	\auto_signaltap_0|acq_data_in_reg [1];
wire	\auto_signaltap_0|acq_data_in_reg[1]~feeder_combout ;
//wire	\auto_signaltap_0|acq_data_in_reg [2];
wire	\auto_signaltap_0|acq_data_in_reg[2]~feeder_combout ;
//wire	\auto_signaltap_0|acq_data_in_reg [3];
//wire	\auto_signaltap_0|acq_data_in_reg [4];
wire	\auto_signaltap_0|acq_data_in_reg[4]~feeder_combout ;
//wire	\auto_signaltap_0|acq_data_in_reg [5];
//wire	\auto_signaltap_0|acq_data_in_reg [6];
wire	\auto_signaltap_0|acq_data_in_reg[6]~feeder_combout ;
//wire	\auto_signaltap_0|acq_data_in_reg [7];
wire	\auto_signaltap_0|acq_data_in_reg[7]~feeder_combout ;
wire	[7:0] \auto_signaltap_0|acq_trigger_in_reg ;
//wire	\auto_signaltap_0|acq_trigger_in_reg [0];
//wire	\auto_signaltap_0|acq_trigger_in_reg [1];
//wire	\auto_signaltap_0|acq_trigger_in_reg [2];
//wire	\auto_signaltap_0|acq_trigger_in_reg [3];
//wire	\auto_signaltap_0|acq_trigger_in_reg [4];
//wire	\auto_signaltap_0|acq_trigger_in_reg [5];
//wire	\auto_signaltap_0|acq_trigger_in_reg [6];
//wire	\auto_signaltap_0|acq_trigger_in_reg [7];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~3_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~5_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~7_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~8_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7]~q ;
wire	[6:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [0];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[0]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [1];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[1]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [2];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[2]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [3];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [4];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[4]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [5];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[5]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [6];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[6]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout ;
wire	[3:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [0];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[0]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [1];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[1]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [2];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[2]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [3];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|Add0~0_combout ;
wire	[3:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [2];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [3];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~10_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~11_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~3_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~5_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~7_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~8_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~9_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal~combout ;
wire	[3:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [3];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter~11_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter~7_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter~8_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter~9_combout ;
wire	[0:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed [0];
wire	[23:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [0];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[0]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [10];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[10]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [11];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[11]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [12];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[12]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [13];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[13]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [14];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[14]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [15];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[15]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [16];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [17];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[17]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [18];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[18]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [19];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[19]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [1];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[1]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [20];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [21];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [22];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [23];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[23]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [2];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[2]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [3];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [5];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[5]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [6];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[6]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [7];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[7]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [8];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[8]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [9];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[9]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|p_match_out~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|p_match_out~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|p_match_out~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|p_match_out~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|p_match_out~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|p_match_out~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|p_match_out~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|p_match_out~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|p_match_out~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|p_match_out~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|p_match_out~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|p_match_out~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|p_match_out~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|p_match_out~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|p_match_out~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|p_match_out~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~q ;
wire	[9:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [1];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[1]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [3];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[3]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [5];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [6];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[6]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [7];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[7]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [8];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[8]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [9];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run~q ;
wire	[3:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [0];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[0]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [1];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[1]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [3];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[3]~feeder_combout ;
wire	[6:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [1];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[1]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [3];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[3]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [5];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[5]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [6];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[6]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X11_Y14_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y14_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y18_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X13_Y18_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y18_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y19_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X18_Y19_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y18_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X22_Y19_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X23_Y19_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ;
wire	[6:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [1];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[1]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [2];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[2]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [3];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[3]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [4];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[4]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [5];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[5]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [6];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[6]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~1 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~10_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~11 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~12_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~3 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~5 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~7 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~8_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~9 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~1 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~10_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~11_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~12 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~13_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~14_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~15 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~16_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~17_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~18 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~19_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~20_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~22_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~3 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~5_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~6 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~7_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~8_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~9 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~3_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|base_address~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|collecting_post_data_var~0_combout ;
wire	[7:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [3];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [5];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [6];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [7];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter~5_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~2_combout ;
wire	[6:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [0];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [1];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[1]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [2];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[2]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [3];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[3]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [4];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[4]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [5];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[5]~feeder_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [6];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[6]~feeder_combout ;
wire	[7:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [0];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[0]~21_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [1];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1]~7_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1]~8 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [2];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2]~10 ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2]~9_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [3];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3]~11_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3]~12 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [4];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4]~13_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4]~14 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [5];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5]~15_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5]~16 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [6];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6]~17_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6]~18 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [7];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[7]~19_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~3_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~5_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~10_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~11_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~12_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~13_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~14_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~15_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~16_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~17_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~3_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~5_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~7_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~8_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~9_combout ;
wire	[16:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [10];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [11];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [12];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [13];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [14];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [15];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [16];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [3];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [5];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [6];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [7];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [8];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [9];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~combout__SyncLoad_X16_Y17_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_comb_bita0~COUT ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_comb_bita0~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_comb_bita1~COUT ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_comb_bita1~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_comb_bita2~combout ;
wire	[2:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [2];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~10_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~11_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~12_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~13_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~14_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~3_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~5_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~7_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~8_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~9_combout ;
wire	[14:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [10];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [11];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [12];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [13];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [14];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [3];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [5];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [6];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [7];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [8];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [9];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena~combout__SyncLoad_X18_Y18_INV ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~3_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~5_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~7_combout ;
wire	[7:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [3];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [5];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [6];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [7];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita0~COUT ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita0~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita1~COUT ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita1~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita2~COUT ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita2~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita3~COUT ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita3~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita4~COUT ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita4~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita5~COUT ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita5~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita6~combout ;
wire	[6:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [3];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [5];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [6];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita0~COUT ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita0~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita1~COUT ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita1~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita2~COUT ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita2~combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~COUT ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~combout ;
wire	[3:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [3];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0_combout__SyncLoad_X17_Y20_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~10_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~11_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~12_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~13_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~14_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~3_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~5_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~7_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~8_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~9_combout ;
wire	[14:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [10];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [11];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [12];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [13];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [14];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [3];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [5];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [6];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [7];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [8];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [9];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~COUT ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~combout ;
wire	[0:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit [0];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0_combout__SyncLoad_X18_Y20_SIG ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9]~feeder_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9]~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[0]~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[10]~10_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[11]~11_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[12]~12_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[13]~13_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[14]~14_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[1]~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[2]~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[3]~3_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[4]~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[5]~5_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[6]~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[7]~7_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[8]~8_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[9]~9_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout ;
wire	[14:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [10];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [11];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [12];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [13];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [14];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [3];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [5];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [6];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [7];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [8];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [9];
wire	[0:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr[0]~feeder_combout ;
wire	[35:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [0];
wire	[17:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [10];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [10];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [11];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [11];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [12];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [12];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [13];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [13];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [14];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [14];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [15];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [15];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [16];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [16];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [17];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [17];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [18];
wire	[17:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [19];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [20];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [21];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [3];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [22];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [23];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [5];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [24];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [6];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [25];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [7];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [26];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [8];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [27];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [9];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [28];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [10];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [29];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [11];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [30];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [12];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [31];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [13];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [32];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [14];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [33];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [15];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [34];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [16];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [35];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [17];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [3];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [3];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [5];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [5];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [6];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [6];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [7];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [7];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [8];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [8];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0_PORTBDATAOUT_bus [9];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [9];
wire	[15:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [0];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [10];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [11];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [12];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [13];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [14];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [15];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [3];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [5];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [6];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [7];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [8];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [9];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~10_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~11_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~12_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~13_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~3_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~5_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~7_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~8_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~9_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ;
wire	[31:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [0];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0]~32_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0]~33 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [10];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~34_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~54_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~55 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [11];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11]~56_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11]~57 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [12];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12]~58_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12]~59 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [13];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13]~60_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13]~61 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [14];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14]~62_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14]~63 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [15];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15]~64_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15]~65 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [16];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16]~66_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16]~67 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [17];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17]~68_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17]~69 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [18];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18]~70_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18]~71 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [19];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19]~72_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19]~73 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [1];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1]~36_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1]~37 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [20];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20]~74_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20]~75 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [21];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21]~76_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21]~77 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [22];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22]~78_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22]~79 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [23];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23]~80_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23]~81 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [24];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24]~82_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24]~83 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [25];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25]~84_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25]~85 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [26];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26]~86_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26]~87 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [27];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27]~88_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27]~89 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [28];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28]~90_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28]~91 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [29];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29]~92_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29]~93 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [2];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2]~38_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2]~39 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [30];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30]~94_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30]~95 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [31];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[31]~96_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [3];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3]~40_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3]~41 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [4];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4]~42_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4]~43 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [5];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5]~44_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5]~45 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [6];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6]~46_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6]~47 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [7];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7]~48_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7]~49 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [8];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8]~50_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8]~51 ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [9];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9]~52_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9]~53 ;
wire	[15:0] \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [0];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout ;
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [10];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [11];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [12];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [13];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [14];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [15];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [1];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [2];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [3];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [4];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [5];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [6];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [7];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [8];
//wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [9];
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~10_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~11_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~12_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~13_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~14_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~15_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~16_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~3_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~5_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~7_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~8_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~9_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~1_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~3_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~4_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~5_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~6_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff~0_combout ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff~q ;
wire	\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout ;
wire	\auto_signaltap_0|~GND~combout ;
wire	\cam_data[0]~input_o ;
wire	\cam_data[1]~input_o ;
wire	\cam_data[2]~input_o ;
wire	\cam_data[3]~input_o ;
wire	\cam_data[4]~input_o ;
wire	\cam_data[5]~input_o ;
wire	\cam_data[6]~input_o ;
wire	\cam_data[7]~input_o ;
wire	\cam_hsync~input_o ;
wire	\cam_pclk~input_o ;
wire	\cam_pclk~input_o_X10_Y9_SIG_VCC ;
wire	\cam_pclk~input_o_X11_Y9_SIG_VCC ;
wire	\cam_pclk~input_o_X13_Y9_SIG_VCC ;
wire	\cam_pclk~input_o_X14_Y8_SIG_VCC ;
wire	\cam_pclk~input_o_X14_Y9_SIG_VCC ;
wire	\cam_pclk~input_o_X16_Y9_SIG_VCC ;
wire	\cam_pclk~input_o_X17_Y9_SIG_VCC ;
wire	\cam_pclk~input_o_X1_Y7_SIG_VCC ;
wire	\cam_pclk~input_o_X2_Y7_SIG_VCC ;
wire	\cam_pclk~input_o_X9_Y7_SIG_VCC ;
wire	\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ;
wire	\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X12_Y9_SIG_SIG ;
wire	\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X13_Y9_SIG_SIG ;
wire	\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X12_Y9_SIG_SIG ;
wire	\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X13_Y7_SIG_SIG ;
wire	\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y9_SIG_SIG ;
wire	\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y9_SIG_SIG ;
wire	\cam_sda~input_o ;
wire	\cam_vsync~input_o ;
wire	\camera_if_inst|Equal0~0_combout ;
wire	\camera_if_inst|Equal0~1_combout ;
wire	\camera_if_inst|Equal0~2_combout ;
wire	\camera_if_inst|Equal0~3_combout ;
wire	\camera_if_inst|Equal0~4_combout ;
wire	\camera_if_inst|Equal1~0_combout ;
wire	\camera_if_inst|Equal1~1_combout ;
wire	\camera_if_inst|Equal2~0_combout ;
wire	\camera_if_inst|Equal3~0_combout ;
wire	\camera_if_inst|Equal3~1_combout ;
wire	\camera_if_inst|Equal3~2_combout ;
wire	\camera_if_inst|Equal3~3_combout ;
wire	\camera_if_inst|Equal3~4_combout ;
wire	\camera_if_inst|Equal4~0_combout ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y9_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y10_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y7_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y11_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y9_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y8_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ;
wire	\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ;
wire	[7:0] \camera_if_inst|cam_data_r0 ;
//wire	\camera_if_inst|cam_data_r0 [0];
//wire	\camera_if_inst|cam_data_r0 [1];
//wire	\camera_if_inst|cam_data_r0 [2];
//wire	\camera_if_inst|cam_data_r0 [3];
//wire	\camera_if_inst|cam_data_r0 [4];
wire	\camera_if_inst|cam_data_r0[4]~feeder_combout ;
//wire	\camera_if_inst|cam_data_r0 [5];
//wire	\camera_if_inst|cam_data_r0 [6];
//wire	\camera_if_inst|cam_data_r0 [7];
wire	[7:0] \camera_if_inst|cam_data_r1 ;
//wire	\camera_if_inst|cam_data_r1 [0];
//wire	\camera_if_inst|cam_data_r1 [1];
//wire	\camera_if_inst|cam_data_r1 [2];
//wire	\camera_if_inst|cam_data_r1 [3];
//wire	\camera_if_inst|cam_data_r1 [4];
//wire	\camera_if_inst|cam_data_r1 [5];
//wire	\camera_if_inst|cam_data_r1 [6];
//wire	\camera_if_inst|cam_data_r1 [7];
wire	\camera_if_inst|cam_data_r1~0_combout ;
wire	\camera_if_inst|cam_data_r1~1_combout ;
wire	\camera_if_inst|cam_data_r1~2_combout ;
wire	\camera_if_inst|cam_data_r1~3_combout ;
wire	\camera_if_inst|cam_data_r1~4_combout ;
wire	\camera_if_inst|cam_data_r1~5_combout ;
wire	\camera_if_inst|cam_data_r1~6_combout ;
wire	\camera_if_inst|cam_data_r1~7_combout ;
wire	[4:0] \camera_if_inst|cam_hsync_r ;
//wire	\camera_if_inst|cam_hsync_r [0];
wire	\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ;
//wire	\camera_if_inst|cam_hsync_r [1];
//wire	\camera_if_inst|cam_hsync_r [2];
//wire	\camera_if_inst|cam_hsync_r [3];
//wire	\camera_if_inst|cam_hsync_r [4];
wire	\camera_if_inst|cam_hsync_r~0_combout ;
wire	\camera_if_inst|cam_hsync_r~1_combout ;
wire	[4:0] \camera_if_inst|cam_vsync_r ;
//wire	\camera_if_inst|cam_vsync_r [0];
wire	\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ;
//wire	\camera_if_inst|cam_vsync_r [1];
//wire	\camera_if_inst|cam_vsync_r [2];
//wire	\camera_if_inst|cam_vsync_r [3];
//wire	\camera_if_inst|cam_vsync_r [4];
wire	[3:0] \camera_if_inst|f_cnt ;
//wire	\camera_if_inst|f_cnt [0];
wire	\camera_if_inst|f_cnt[0]~5_combout ;
//wire	\camera_if_inst|f_cnt [1];
wire	\camera_if_inst|f_cnt[1]~4_combout ;
//wire	\camera_if_inst|f_cnt [2];
wire	\camera_if_inst|f_cnt[2]~3_combout ;
//wire	\camera_if_inst|f_cnt [3];
wire	\camera_if_inst|f_cnt[3]~2_combout ;
wire	\camera_if_inst|f_cnt[3]~6_combout ;
wire	[15:0] \camera_if_inst|h_cnt ;
//wire	\camera_if_inst|h_cnt [0];
wire	\camera_if_inst|h_cnt[0]~16_combout ;
wire	\camera_if_inst|h_cnt[0]~17 ;
//wire	\camera_if_inst|h_cnt [10];
wire	\camera_if_inst|h_cnt[10]~36_combout ;
wire	\camera_if_inst|h_cnt[10]~37 ;
//wire	\camera_if_inst|h_cnt [11];
wire	\camera_if_inst|h_cnt[11]~38_combout ;
wire	\camera_if_inst|h_cnt[11]~39 ;
//wire	\camera_if_inst|h_cnt [12];
wire	\camera_if_inst|h_cnt[12]~40_combout ;
wire	\camera_if_inst|h_cnt[12]~41 ;
//wire	\camera_if_inst|h_cnt [13];
wire	\camera_if_inst|h_cnt[13]~42_combout ;
wire	\camera_if_inst|h_cnt[13]~43 ;
//wire	\camera_if_inst|h_cnt [14];
wire	\camera_if_inst|h_cnt[14]~44_combout ;
wire	\camera_if_inst|h_cnt[14]~45 ;
//wire	\camera_if_inst|h_cnt [15];
wire	\camera_if_inst|h_cnt[15]~46_combout ;
//wire	\camera_if_inst|h_cnt [1];
wire	\camera_if_inst|h_cnt[1]~18_combout ;
wire	\camera_if_inst|h_cnt[1]~19 ;
//wire	\camera_if_inst|h_cnt [2];
wire	\camera_if_inst|h_cnt[2]~20_combout ;
wire	\camera_if_inst|h_cnt[2]~21 ;
//wire	\camera_if_inst|h_cnt [3];
wire	\camera_if_inst|h_cnt[3]~22_combout ;
wire	\camera_if_inst|h_cnt[3]~23 ;
//wire	\camera_if_inst|h_cnt [4];
wire	\camera_if_inst|h_cnt[4]~24_combout ;
wire	\camera_if_inst|h_cnt[4]~25 ;
//wire	\camera_if_inst|h_cnt [5];
wire	\camera_if_inst|h_cnt[5]~26_combout ;
wire	\camera_if_inst|h_cnt[5]~27 ;
//wire	\camera_if_inst|h_cnt [6];
wire	\camera_if_inst|h_cnt[6]~28_combout ;
wire	\camera_if_inst|h_cnt[6]~29 ;
//wire	\camera_if_inst|h_cnt [7];
wire	\camera_if_inst|h_cnt[7]~30_combout ;
wire	\camera_if_inst|h_cnt[7]~31 ;
//wire	\camera_if_inst|h_cnt [8];
wire	\camera_if_inst|h_cnt[8]~32_combout ;
wire	\camera_if_inst|h_cnt[8]~33 ;
//wire	\camera_if_inst|h_cnt [9];
wire	\camera_if_inst|h_cnt[9]~34_combout ;
wire	\camera_if_inst|h_cnt[9]~35 ;
wire	[7:0] \camera_if_inst|u_I2C_AV_Config|LUT_INDEX ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0]~22_combout ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1]~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1]~8 ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2]~10 ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2]~9_combout ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3]~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3]~12 ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4]~14_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4]~15 ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5]~16_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5]~17 ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6]~18_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6]~19 ;
//wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7];
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~20_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan0~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan0~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan0~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan0~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan1~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|Selector3~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|Selector3~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|Selector3~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~feeder_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~q ;
wire	\camera_if_inst|u_I2C_AV_Config|i2c_en_r1~q ;
wire	\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ;
wire	[15:0] \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [0];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0]~16_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0]~17 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [10];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10]~36_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10]~37 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [11];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11]~38_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11]~39 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [12];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12]~40_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12]~41 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [13];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13]~42_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13]~43 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [14];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14]~44_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14]~45 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [15];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15]~46_combout ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [1];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1]~18_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1]~19 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [2];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2]~20_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2]~21 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [3];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3]~22_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3]~23 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [4];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4]~24_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4]~25 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [5];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5]~26_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5]~27 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [6];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6]~28_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6]~29 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [7];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7]~30_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7]~31 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [8];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8]~32_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8]~33 ;
//wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [9];
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9]~34_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9]~35 ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~q ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X19_Y8_INV ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_GO~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_WR~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST.00~q ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST.10~q ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST~12_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|mSetup_ST~13_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACK~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACK~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|ACK~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|END~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Equal0~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Equal0~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Equal3~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Equal3~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Equal5~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~12_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~13_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~14_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~15_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~16_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~17_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~18_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~19_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~20_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~21_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~22_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~23_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~24_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~25_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~26_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~27_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~28_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~29_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~30_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~31_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Mux1~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SDO~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SDO~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SDO~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SDO~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SDO~4_combout ;
wire	[5:0] \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER ;
//wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0];
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0]~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0]~7 ;
//wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1];
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1]~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1]~9 ;
//wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2];
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2]~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2]~11 ;
//wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3];
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3]~13_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3]~14 ;
//wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4];
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4]~15_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4]~16 ;
//wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5];
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~17_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector2~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector6~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector8~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector9~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|Selector9~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|comb~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u0|comb~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8_combout ;
wire	\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9_combout ;
wire	[15:0] \camera_if_inst|v_cnt ;
//wire	\camera_if_inst|v_cnt [0];
wire	\camera_if_inst|v_cnt[0]~16_combout ;
wire	\camera_if_inst|v_cnt[0]~17 ;
//wire	\camera_if_inst|v_cnt [10];
wire	\camera_if_inst|v_cnt[10]~18_combout ;
wire	\camera_if_inst|v_cnt[10]~37_combout ;
wire	\camera_if_inst|v_cnt[10]~38 ;
//wire	\camera_if_inst|v_cnt [11];
wire	\camera_if_inst|v_cnt[11]~39_combout ;
wire	\camera_if_inst|v_cnt[11]~40 ;
//wire	\camera_if_inst|v_cnt [12];
wire	\camera_if_inst|v_cnt[12]~41_combout ;
wire	\camera_if_inst|v_cnt[12]~42 ;
//wire	\camera_if_inst|v_cnt [13];
wire	\camera_if_inst|v_cnt[13]~43_combout ;
wire	\camera_if_inst|v_cnt[13]~44 ;
//wire	\camera_if_inst|v_cnt [14];
wire	\camera_if_inst|v_cnt[14]~45_combout ;
wire	\camera_if_inst|v_cnt[14]~46 ;
//wire	\camera_if_inst|v_cnt [15];
wire	\camera_if_inst|v_cnt[15]~47_combout ;
//wire	\camera_if_inst|v_cnt [1];
wire	\camera_if_inst|v_cnt[1]~19_combout ;
wire	\camera_if_inst|v_cnt[1]~20 ;
//wire	\camera_if_inst|v_cnt [2];
wire	\camera_if_inst|v_cnt[2]~21_combout ;
wire	\camera_if_inst|v_cnt[2]~22 ;
//wire	\camera_if_inst|v_cnt [3];
wire	\camera_if_inst|v_cnt[3]~23_combout ;
wire	\camera_if_inst|v_cnt[3]~24 ;
//wire	\camera_if_inst|v_cnt [4];
wire	\camera_if_inst|v_cnt[4]~25_combout ;
wire	\camera_if_inst|v_cnt[4]~26 ;
//wire	\camera_if_inst|v_cnt [5];
wire	\camera_if_inst|v_cnt[5]~27_combout ;
wire	\camera_if_inst|v_cnt[5]~28 ;
//wire	\camera_if_inst|v_cnt [6];
wire	\camera_if_inst|v_cnt[6]~29_combout ;
wire	\camera_if_inst|v_cnt[6]~30 ;
//wire	\camera_if_inst|v_cnt [7];
wire	\camera_if_inst|v_cnt[7]~31_combout ;
wire	\camera_if_inst|v_cnt[7]~32 ;
//wire	\camera_if_inst|v_cnt [8];
wire	\camera_if_inst|v_cnt[8]~33_combout ;
wire	\camera_if_inst|v_cnt[8]~34 ;
//wire	\camera_if_inst|v_cnt [9];
wire	\camera_if_inst|v_cnt[9]~35_combout ;
wire	\camera_if_inst|v_cnt[9]~36 ;
wire	\clk_25m~0_combout ;
wire	\clk_25m~clkctrl_outclk ;
wire	\clk_25m~clkctrl_outclk_X10_Y9_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X11_Y9_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X13_Y10_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X14_Y10_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X14_Y11_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X16_Y8_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X17_Y9_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X23_Y16_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X24_Y12_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X24_Y16_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X25_Y12_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk_X25_Y15_SIG_VCC ;
wire	\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X13_Y10_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X13_Y7_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y10_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y8_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y12_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y13_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y12_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y13_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y14_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y15_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[4]~13_combout_X24_Y15_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X26_Y16_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout_X25_Y13_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y14_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y15_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X25_Y15_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y16_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X24_Y16_SIG_SIG ;
wire	\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X26_Y16_SIG_SIG ;
wire	\clk_25m~q ;
wire	\clk~input_o ;
wire	\clk~inputclkctrl_outclk ;
wire	\clk~inputclkctrl_outclk_X11_Y14_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X11_Y16_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X12_Y18_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X13_Y16_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X13_Y18_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X14_Y14_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X14_Y16_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X14_Y18_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X16_Y16_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X18_Y19_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X21_Y18_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X21_Y20_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X24_Y18_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ;
wire	\clk~inputclkctrl_outclk_X33_Y12_SIG_VCC ;
wire	\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X16_Y14_SIG_SIG ;
wire	\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X22_Y19_SIG_SIG ;
wire	\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X23_Y19_SIG_SIG ;
wire	\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X16_Y14_SIG_SIG ;
wire	\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X22_Y19_SIG_SIG ;
wire	\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X24_Y19_SIG_SIG ;
wire	\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0_combout_X17_Y14_SIG_SIG ;
wire	\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y18_SIG_SIG ;
wire	\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y19_SIG_SIG ;
wire	\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y18_SIG_SIG ;
wire	\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y19_SIG_SIG ;
wire	\clk~inputclkctrl_outclk__reset_init[5]_X33_Y12_SIG_INV ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita0~COUT ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita0~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~COUT ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~combout ;
wire	[1:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [1];
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [0];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [10];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [2];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [3];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [4];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [5];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9]~feeder_combout ;
wire	[31:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [18];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [19];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [20];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [21];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [22];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [23];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [24];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [25];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [26];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [27];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [28];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [29];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [30];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [31];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|q_b [9];
wire	[7:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [0];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [9];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0_PORTBDATAOUT_bus [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [16];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [9];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [8];
wire	[7:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [0];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [9];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1_PORTBDATAOUT_bus [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [16];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [9];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [8];
wire	[7:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [0];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [9];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2_PORTBDATAOUT_bus [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [16];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [9];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [8];
wire	[7:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6_PORTBDATAOUT_bus ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6_PORTBDATAOUT_bus [0];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [9];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6_PORTBDATAOUT_bus [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6_PORTBDATAOUT_bus [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6_PORTBDATAOUT_bus [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6_PORTBDATAOUT_bus [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6_PORTBDATAOUT_bus [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6_PORTBDATAOUT_bus [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6_PORTBDATAOUT_bus [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [16];
wire	[17:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [12];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [13];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [14];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [15];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [16];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [9];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [17];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [8];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11_cout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~13 ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~15 ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~17 ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1_cout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3_cout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5_cout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7_cout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9_cout ;
wire	[11:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~1_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~2_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~3_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~5_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|data_wire[2]~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~10_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~1_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~7_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~8_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~9_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ;
wire	[2:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [2];
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [0];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0]~0_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [1];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9]~feeder_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor0~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor1~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor2~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor3~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor4~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor5~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor6~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor7~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor8~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor9~combout ;
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [9];
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor0~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor1~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor2~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor3~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor4~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor5~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor6~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor7~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor8~combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor9~combout ;
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [10];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [1];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [2];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [3];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [6];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [7];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9]~feeder_combout ;
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [7];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9]~feeder_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~1_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~2_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~3_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~5_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|data_wire[2]~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~10_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~6_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~7_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~8_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~9_combout ;
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [10];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10]~0_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1]~8_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2]~7_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3]~9_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4]~5_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5]~6_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6]~3_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7]~4_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8]~1_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9]~2_combout ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1~q ;
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2~q ;
wire	[12:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0]~0_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [11];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [12];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9]~feeder_combout ;
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [0];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [10];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [1];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [2];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [3];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [4];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [5];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [6];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [7];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9]~feeder_combout ;
wire	[10:0] \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [0];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [10];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [1];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [2];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [3];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [4];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [5];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [6];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [7];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7]~feeder_combout ;
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [8];
//wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [9];
wire	\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9]~feeder_combout ;
wire	[31:0] \cmos1_fifo_inst|q ;
//wire	\cmos1_fifo_inst|q [0];
//wire	\cmos1_fifo_inst|q [10];
//wire	\cmos1_fifo_inst|q [11];
//wire	\cmos1_fifo_inst|q [12];
//wire	\cmos1_fifo_inst|q [13];
//wire	\cmos1_fifo_inst|q [14];
//wire	\cmos1_fifo_inst|q [15];
//wire	\cmos1_fifo_inst|q [16];
//wire	\cmos1_fifo_inst|q [17];
//wire	\cmos1_fifo_inst|q [18];
//wire	\cmos1_fifo_inst|q [19];
//wire	\cmos1_fifo_inst|q [1];
//wire	\cmos1_fifo_inst|q [20];
//wire	\cmos1_fifo_inst|q [21];
//wire	\cmos1_fifo_inst|q [22];
//wire	\cmos1_fifo_inst|q [23];
//wire	\cmos1_fifo_inst|q [24];
//wire	\cmos1_fifo_inst|q [25];
//wire	\cmos1_fifo_inst|q [26];
//wire	\cmos1_fifo_inst|q [27];
//wire	\cmos1_fifo_inst|q [28];
//wire	\cmos1_fifo_inst|q [29];
//wire	\cmos1_fifo_inst|q [2];
//wire	\cmos1_fifo_inst|q [30];
//wire	\cmos1_fifo_inst|q [31];
//wire	\cmos1_fifo_inst|q [3];
//wire	\cmos1_fifo_inst|q [4];
//wire	\cmos1_fifo_inst|q [5];
//wire	\cmos1_fifo_inst|q [6];
//wire	\cmos1_fifo_inst|q [7];
//wire	\cmos1_fifo_inst|q [8];
//wire	\cmos1_fifo_inst|q [9];
wire	\cmos1_fifo_inst|q~0_combout ;
wire	\cmos1_fifo_inst|q~10_combout ;
wire	\cmos1_fifo_inst|q~11_combout ;
wire	\cmos1_fifo_inst|q~12_combout ;
wire	\cmos1_fifo_inst|q~13_combout ;
wire	\cmos1_fifo_inst|q~14_combout ;
wire	\cmos1_fifo_inst|q~15_combout ;
wire	\cmos1_fifo_inst|q~16_combout ;
wire	\cmos1_fifo_inst|q~17_combout ;
wire	\cmos1_fifo_inst|q~18_combout ;
wire	\cmos1_fifo_inst|q~19_combout ;
wire	\cmos1_fifo_inst|q~1_combout ;
wire	\cmos1_fifo_inst|q~20_combout ;
wire	\cmos1_fifo_inst|q~21_combout ;
wire	\cmos1_fifo_inst|q~22_combout ;
wire	\cmos1_fifo_inst|q~23_combout ;
wire	\cmos1_fifo_inst|q~24_combout ;
wire	\cmos1_fifo_inst|q~25_combout ;
wire	\cmos1_fifo_inst|q~26_combout ;
wire	\cmos1_fifo_inst|q~27_combout ;
wire	\cmos1_fifo_inst|q~28_combout ;
wire	\cmos1_fifo_inst|q~29_combout ;
wire	\cmos1_fifo_inst|q~2_combout ;
wire	\cmos1_fifo_inst|q~30_combout ;
wire	\cmos1_fifo_inst|q~31_combout ;
wire	\cmos1_fifo_inst|q~3_combout ;
wire	\cmos1_fifo_inst|q~4_combout ;
wire	\cmos1_fifo_inst|q~5_combout ;
wire	\cmos1_fifo_inst|q~6_combout ;
wire	\cmos1_fifo_inst|q~7_combout ;
wire	\cmos1_fifo_inst|q~8_combout ;
wire	\cmos1_fifo_inst|q~9_combout ;
tri1	devclrn;
tri1	devoe;
tri1	devpor;
wire	\e_rx[0]~input_o ;
wire	\e_rx[1]~input_o ;
wire	\e_rxclk~input_o ;
wire	\e_rxclk~input_o_X33_Y16_INV_VCC ;
wire	\e_rxclk~input_o__mii_to_rmii_inst|tx_dv_reg~q_X33_Y16_SIG_SIG ;
wire	\e_rxdv~input_o ;
wire	\e_rxer~input_o ;
wire	[31:0] \eth_udp_inst|crc32_inst|crc_data ;
//wire	\eth_udp_inst|crc32_inst|crc_data [0];
//wire	\eth_udp_inst|crc32_inst|crc_data [10];
//wire	\eth_udp_inst|crc32_inst|crc_data [11];
//wire	\eth_udp_inst|crc32_inst|crc_data [12];
//wire	\eth_udp_inst|crc32_inst|crc_data [13];
//wire	\eth_udp_inst|crc32_inst|crc_data [14];
//wire	\eth_udp_inst|crc32_inst|crc_data [15];
//wire	\eth_udp_inst|crc32_inst|crc_data [16];
//wire	\eth_udp_inst|crc32_inst|crc_data [17];
//wire	\eth_udp_inst|crc32_inst|crc_data [18];
//wire	\eth_udp_inst|crc32_inst|crc_data [19];
//wire	\eth_udp_inst|crc32_inst|crc_data [1];
//wire	\eth_udp_inst|crc32_inst|crc_data [20];
//wire	\eth_udp_inst|crc32_inst|crc_data [21];
//wire	\eth_udp_inst|crc32_inst|crc_data [22];
//wire	\eth_udp_inst|crc32_inst|crc_data [23];
//wire	\eth_udp_inst|crc32_inst|crc_data [24];
//wire	\eth_udp_inst|crc32_inst|crc_data [25];
//wire	\eth_udp_inst|crc32_inst|crc_data [26];
//wire	\eth_udp_inst|crc32_inst|crc_data [27];
//wire	\eth_udp_inst|crc32_inst|crc_data [28];
//wire	\eth_udp_inst|crc32_inst|crc_data [29];
wire	\eth_udp_inst|crc32_inst|crc_data[29]~9_combout ;
//wire	\eth_udp_inst|crc32_inst|crc_data [2];
//wire	\eth_udp_inst|crc32_inst|crc_data [30];
//wire	\eth_udp_inst|crc32_inst|crc_data [31];
//wire	\eth_udp_inst|crc32_inst|crc_data [3];
//wire	\eth_udp_inst|crc32_inst|crc_data [4];
//wire	\eth_udp_inst|crc32_inst|crc_data [5];
//wire	\eth_udp_inst|crc32_inst|crc_data [6];
//wire	\eth_udp_inst|crc32_inst|crc_data [7];
//wire	\eth_udp_inst|crc32_inst|crc_data [8];
//wire	\eth_udp_inst|crc32_inst|crc_data [9];
wire	\eth_udp_inst|crc32_inst|crc_data~10_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~11_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~12_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~13_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~14_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~15_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~16_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~17_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~18_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~19_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~20_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~21_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~22_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~23_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~24_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~25_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~26_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~27_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~28_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~29_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~30_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~31_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~32_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~33_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~34_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~35_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~36_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~37_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~38_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~39_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~40_combout ;
wire	\eth_udp_inst|crc32_inst|crc_data~8_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next[28]~1_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next[29]~0_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next~2_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next~3_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next~4_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next~5_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next~6_combout ;
wire	\eth_udp_inst|crc32_inst|crc_next~7_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~1 ;
wire	\eth_udp_inst|ip_send_inst|Add13~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~11 ;
wire	\eth_udp_inst|ip_send_inst|Add13~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~13 ;
wire	\eth_udp_inst|ip_send_inst|Add13~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~15 ;
wire	\eth_udp_inst|ip_send_inst|Add13~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~17 ;
wire	\eth_udp_inst|ip_send_inst|Add13~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~19 ;
wire	\eth_udp_inst|ip_send_inst|Add13~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~21 ;
wire	\eth_udp_inst|ip_send_inst|Add13~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~23 ;
wire	\eth_udp_inst|ip_send_inst|Add13~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~25 ;
wire	\eth_udp_inst|ip_send_inst|Add13~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~27 ;
wire	\eth_udp_inst|ip_send_inst|Add13~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~29 ;
wire	\eth_udp_inst|ip_send_inst|Add13~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~3 ;
wire	\eth_udp_inst|ip_send_inst|Add13~30_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~5 ;
wire	\eth_udp_inst|ip_send_inst|Add13~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~7 ;
wire	\eth_udp_inst|ip_send_inst|Add13~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add13~9 ;
wire	\eth_udp_inst|ip_send_inst|Add2~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~1 ;
wire	\eth_udp_inst|ip_send_inst|Add2~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~11 ;
wire	\eth_udp_inst|ip_send_inst|Add2~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~13 ;
wire	\eth_udp_inst|ip_send_inst|Add2~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~15 ;
wire	\eth_udp_inst|ip_send_inst|Add2~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~17 ;
wire	\eth_udp_inst|ip_send_inst|Add2~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~19 ;
wire	\eth_udp_inst|ip_send_inst|Add2~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~21 ;
wire	\eth_udp_inst|ip_send_inst|Add2~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~23 ;
wire	\eth_udp_inst|ip_send_inst|Add2~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~25 ;
wire	\eth_udp_inst|ip_send_inst|Add2~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~27 ;
wire	\eth_udp_inst|ip_send_inst|Add2~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~3 ;
wire	\eth_udp_inst|ip_send_inst|Add2~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~5 ;
wire	\eth_udp_inst|ip_send_inst|Add2~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~7 ;
wire	\eth_udp_inst|ip_send_inst|Add2~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add2~9 ;
wire	\eth_udp_inst|ip_send_inst|Add3~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add3~1 ;
wire	\eth_udp_inst|ip_send_inst|Add3~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add3~3 ;
wire	\eth_udp_inst|ip_send_inst|Add3~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~1 ;
wire	\eth_udp_inst|ip_send_inst|Add4~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~11 ;
wire	\eth_udp_inst|ip_send_inst|Add4~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~13 ;
wire	\eth_udp_inst|ip_send_inst|Add4~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~15 ;
wire	\eth_udp_inst|ip_send_inst|Add4~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~17 ;
wire	\eth_udp_inst|ip_send_inst|Add4~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~19 ;
wire	\eth_udp_inst|ip_send_inst|Add4~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~21 ;
wire	\eth_udp_inst|ip_send_inst|Add4~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~23 ;
wire	\eth_udp_inst|ip_send_inst|Add4~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~25 ;
wire	\eth_udp_inst|ip_send_inst|Add4~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~27 ;
wire	\eth_udp_inst|ip_send_inst|Add4~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~29 ;
wire	\eth_udp_inst|ip_send_inst|Add4~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~3 ;
wire	\eth_udp_inst|ip_send_inst|Add4~30_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~31 ;
wire	\eth_udp_inst|ip_send_inst|Add4~32_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~33 ;
wire	\eth_udp_inst|ip_send_inst|Add4~34_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~5 ;
wire	\eth_udp_inst|ip_send_inst|Add4~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~7 ;
wire	\eth_udp_inst|ip_send_inst|Add4~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add4~9 ;
wire	\eth_udp_inst|ip_send_inst|Add5~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~1 ;
wire	\eth_udp_inst|ip_send_inst|Add5~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~11 ;
wire	\eth_udp_inst|ip_send_inst|Add5~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~13 ;
wire	\eth_udp_inst|ip_send_inst|Add5~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~15 ;
wire	\eth_udp_inst|ip_send_inst|Add5~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~17 ;
wire	\eth_udp_inst|ip_send_inst|Add5~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~19 ;
wire	\eth_udp_inst|ip_send_inst|Add5~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~21 ;
wire	\eth_udp_inst|ip_send_inst|Add5~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~23 ;
wire	\eth_udp_inst|ip_send_inst|Add5~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~25 ;
wire	\eth_udp_inst|ip_send_inst|Add5~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~27 ;
wire	\eth_udp_inst|ip_send_inst|Add5~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~29 ;
wire	\eth_udp_inst|ip_send_inst|Add5~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~3 ;
wire	\eth_udp_inst|ip_send_inst|Add5~30_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~31 ;
wire	\eth_udp_inst|ip_send_inst|Add5~32_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~33 ;
wire	\eth_udp_inst|ip_send_inst|Add5~34_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~5 ;
wire	\eth_udp_inst|ip_send_inst|Add5~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~7 ;
wire	\eth_udp_inst|ip_send_inst|Add5~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add5~9 ;
wire	\eth_udp_inst|ip_send_inst|Add6~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~1 ;
wire	\eth_udp_inst|ip_send_inst|Add6~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~11 ;
wire	\eth_udp_inst|ip_send_inst|Add6~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~13 ;
wire	\eth_udp_inst|ip_send_inst|Add6~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~15 ;
wire	\eth_udp_inst|ip_send_inst|Add6~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~17 ;
wire	\eth_udp_inst|ip_send_inst|Add6~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~19 ;
wire	\eth_udp_inst|ip_send_inst|Add6~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~21 ;
wire	\eth_udp_inst|ip_send_inst|Add6~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~23 ;
wire	\eth_udp_inst|ip_send_inst|Add6~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~25 ;
wire	\eth_udp_inst|ip_send_inst|Add6~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~27 ;
wire	\eth_udp_inst|ip_send_inst|Add6~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~3 ;
wire	\eth_udp_inst|ip_send_inst|Add6~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~5 ;
wire	\eth_udp_inst|ip_send_inst|Add6~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~7 ;
wire	\eth_udp_inst|ip_send_inst|Add6~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add6~9 ;
wire	\eth_udp_inst|ip_send_inst|Add7~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~1 ;
wire	\eth_udp_inst|ip_send_inst|Add7~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~11 ;
wire	\eth_udp_inst|ip_send_inst|Add7~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~13 ;
wire	\eth_udp_inst|ip_send_inst|Add7~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~15 ;
wire	\eth_udp_inst|ip_send_inst|Add7~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~17 ;
wire	\eth_udp_inst|ip_send_inst|Add7~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~19 ;
wire	\eth_udp_inst|ip_send_inst|Add7~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~21 ;
wire	\eth_udp_inst|ip_send_inst|Add7~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~23 ;
wire	\eth_udp_inst|ip_send_inst|Add7~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~25 ;
wire	\eth_udp_inst|ip_send_inst|Add7~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~27 ;
wire	\eth_udp_inst|ip_send_inst|Add7~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~29 ;
wire	\eth_udp_inst|ip_send_inst|Add7~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~3 ;
wire	\eth_udp_inst|ip_send_inst|Add7~30_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~31 ;
wire	\eth_udp_inst|ip_send_inst|Add7~32_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~5 ;
wire	\eth_udp_inst|ip_send_inst|Add7~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~7 ;
wire	\eth_udp_inst|ip_send_inst|Add7~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add7~9 ;
wire	\eth_udp_inst|ip_send_inst|Add8~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~1 ;
wire	\eth_udp_inst|ip_send_inst|Add8~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~11 ;
wire	\eth_udp_inst|ip_send_inst|Add8~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~13 ;
wire	\eth_udp_inst|ip_send_inst|Add8~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~15 ;
wire	\eth_udp_inst|ip_send_inst|Add8~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~17 ;
wire	\eth_udp_inst|ip_send_inst|Add8~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~19 ;
wire	\eth_udp_inst|ip_send_inst|Add8~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~21 ;
wire	\eth_udp_inst|ip_send_inst|Add8~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~23 ;
wire	\eth_udp_inst|ip_send_inst|Add8~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~25 ;
wire	\eth_udp_inst|ip_send_inst|Add8~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~27 ;
wire	\eth_udp_inst|ip_send_inst|Add8~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~29 ;
wire	\eth_udp_inst|ip_send_inst|Add8~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~3 ;
wire	\eth_udp_inst|ip_send_inst|Add8~30_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~5 ;
wire	\eth_udp_inst|ip_send_inst|Add8~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~7 ;
wire	\eth_udp_inst|ip_send_inst|Add8~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add8~9 ;
wire	\eth_udp_inst|ip_send_inst|Add9~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~1 ;
wire	\eth_udp_inst|ip_send_inst|Add9~10_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~11 ;
wire	\eth_udp_inst|ip_send_inst|Add9~12_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~13 ;
wire	\eth_udp_inst|ip_send_inst|Add9~14_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~15 ;
wire	\eth_udp_inst|ip_send_inst|Add9~16_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~17 ;
wire	\eth_udp_inst|ip_send_inst|Add9~18_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~19 ;
wire	\eth_udp_inst|ip_send_inst|Add9~20_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~21 ;
wire	\eth_udp_inst|ip_send_inst|Add9~22_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~23 ;
wire	\eth_udp_inst|ip_send_inst|Add9~24_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~25 ;
wire	\eth_udp_inst|ip_send_inst|Add9~26_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~27 ;
wire	\eth_udp_inst|ip_send_inst|Add9~28_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~29 ;
wire	\eth_udp_inst|ip_send_inst|Add9~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~3 ;
wire	\eth_udp_inst|ip_send_inst|Add9~30_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~31 ;
wire	\eth_udp_inst|ip_send_inst|Add9~32_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~33 ;
wire	\eth_udp_inst|ip_send_inst|Add9~34_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~35 ;
wire	\eth_udp_inst|ip_send_inst|Add9~36_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~5 ;
wire	\eth_udp_inst|ip_send_inst|Add9~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~7 ;
wire	\eth_udp_inst|ip_send_inst|Add9~8_combout ;
wire	\eth_udp_inst|ip_send_inst|Add9~9 ;
wire	\eth_udp_inst|ip_send_inst|Equal1~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal1~1_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y14_SIG ;
wire	\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y15_SIG ;
wire	\eth_udp_inst|ip_send_inst|Equal8~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal8~1_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal8~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal8~3_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal8~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal8~5_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal8~6_combout ;
wire	\eth_udp_inst|ip_send_inst|Equal9~0_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~0_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~1_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~2_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~3_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~4_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~5_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~6_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan1~7_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan2~0_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan2~1_combout ;
wire	\eth_udp_inst|ip_send_inst|LessThan2~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux13~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux13~1_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux13~2_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux13~3_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux13~4_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux16~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux17~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux17~1_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux20~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux21~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux24~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux24~1_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux25~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux27~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux28~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux29~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux31~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux32~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux33~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux35~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux35~1_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux36~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux37~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux39~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux40~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux41~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux43~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux44~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux45~0_combout ;
wire	\eth_udp_inst|ip_send_inst|Mux47~0_combout ;
wire	\eth_udp_inst|ip_send_inst|always10~0_combout ;
wire	\eth_udp_inst|ip_send_inst|always11~0_combout ;
wire	\eth_udp_inst|ip_send_inst|always13~0_combout ;
wire	\eth_udp_inst|ip_send_inst|always16~0_combout ;
wire	\eth_udp_inst|ip_send_inst|always3~2_combout ;
wire	\eth_udp_inst|ip_send_inst|always3~3_combout ;
wire	\eth_udp_inst|ip_send_inst|always3~4_combout ;
wire	\eth_udp_inst|ip_send_inst|always7~0_combout ;
wire	\eth_udp_inst|ip_send_inst|always7~1_combout ;
wire	[31:0] \eth_udp_inst|ip_send_inst|check_sum ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [0];
wire	\eth_udp_inst|ip_send_inst|check_sum[0]~17_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[0]~18 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [10];
wire	\eth_udp_inst|ip_send_inst|check_sum[10]~37_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[10]~38 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [11];
wire	\eth_udp_inst|ip_send_inst|check_sum[11]~39_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[11]~40 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [12];
wire	\eth_udp_inst|ip_send_inst|check_sum[12]~41_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[12]~42 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [13];
wire	\eth_udp_inst|ip_send_inst|check_sum[13]~43_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[13]~44 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [14];
wire	\eth_udp_inst|ip_send_inst|check_sum[14]~45_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[14]~46 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [15];
wire	\eth_udp_inst|ip_send_inst|check_sum[15]~48_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[15]~49 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [16];
wire	\eth_udp_inst|ip_send_inst|check_sum[16]~52_combout ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [17];
//wire	\eth_udp_inst|ip_send_inst|check_sum [18];
//wire	\eth_udp_inst|ip_send_inst|check_sum [19];
//wire	\eth_udp_inst|ip_send_inst|check_sum [1];
wire	\eth_udp_inst|ip_send_inst|check_sum[1]~19_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[1]~20 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [20];
//wire	\eth_udp_inst|ip_send_inst|check_sum [21];
//wire	\eth_udp_inst|ip_send_inst|check_sum [22];
//wire	\eth_udp_inst|ip_send_inst|check_sum [23];
//wire	\eth_udp_inst|ip_send_inst|check_sum [24];
//wire	\eth_udp_inst|ip_send_inst|check_sum [25];
//wire	\eth_udp_inst|ip_send_inst|check_sum [26];
//wire	\eth_udp_inst|ip_send_inst|check_sum [27];
//wire	\eth_udp_inst|ip_send_inst|check_sum [28];
//wire	\eth_udp_inst|ip_send_inst|check_sum [29];
//wire	\eth_udp_inst|ip_send_inst|check_sum [2];
wire	\eth_udp_inst|ip_send_inst|check_sum[2]~21_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[2]~22 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [30];
//wire	\eth_udp_inst|ip_send_inst|check_sum [31];
//wire	\eth_udp_inst|ip_send_inst|check_sum [3];
wire	\eth_udp_inst|ip_send_inst|check_sum[3]~23_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[3]~24 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [4];
wire	\eth_udp_inst|ip_send_inst|check_sum[4]~25_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[4]~26 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [5];
wire	\eth_udp_inst|ip_send_inst|check_sum[5]~27_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[5]~28 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [6];
wire	\eth_udp_inst|ip_send_inst|check_sum[6]~29_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[6]~30 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [7];
wire	\eth_udp_inst|ip_send_inst|check_sum[7]~31_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[7]~32 ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [8];
wire	\eth_udp_inst|ip_send_inst|check_sum[8]~33_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[8]~34 ;
wire	\eth_udp_inst|ip_send_inst|check_sum[8]~47_combout ;
//wire	\eth_udp_inst|ip_send_inst|check_sum [9];
wire	\eth_udp_inst|ip_send_inst|check_sum[9]~35_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum[9]~36 ;
wire	\eth_udp_inst|ip_send_inst|check_sum~50_combout ;
wire	\eth_udp_inst|ip_send_inst|check_sum~51_combout ;
wire	[4:0] \eth_udp_inst|ip_send_inst|cnt ;
//wire	\eth_udp_inst|ip_send_inst|cnt [0];
wire	\eth_udp_inst|ip_send_inst|cnt[0]~5_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt[0]~6 ;
//wire	\eth_udp_inst|ip_send_inst|cnt [1];
wire	\eth_udp_inst|ip_send_inst|cnt[1]~7_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt[1]~8 ;
//wire	\eth_udp_inst|ip_send_inst|cnt [2];
wire	\eth_udp_inst|ip_send_inst|cnt[2]~10 ;
wire	\eth_udp_inst|ip_send_inst|cnt[2]~9_combout ;
//wire	\eth_udp_inst|ip_send_inst|cnt [3];
wire	\eth_udp_inst|ip_send_inst|cnt[3]~14_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt[3]~15 ;
//wire	\eth_udp_inst|ip_send_inst|cnt [4];
wire	\eth_udp_inst|ip_send_inst|cnt[4]~11_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt[4]~11_combout__SyncReset_X24_Y15_SIG ;
wire	\eth_udp_inst|ip_send_inst|cnt[4]~12_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt[4]~13_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt[4]~16_combout ;
wire	[4:0] \eth_udp_inst|ip_send_inst|cnt_add ;
//wire	\eth_udp_inst|ip_send_inst|cnt_add [0];
wire	\eth_udp_inst|ip_send_inst|cnt_add[0]~5_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_add[0]~6 ;
//wire	\eth_udp_inst|ip_send_inst|cnt_add [1];
wire	\eth_udp_inst|ip_send_inst|cnt_add[1]~7_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_add[1]~8 ;
//wire	\eth_udp_inst|ip_send_inst|cnt_add [2];
wire	\eth_udp_inst|ip_send_inst|cnt_add[2]~10 ;
wire	\eth_udp_inst|ip_send_inst|cnt_add[2]~9_combout ;
//wire	\eth_udp_inst|ip_send_inst|cnt_add [3];
wire	\eth_udp_inst|ip_send_inst|cnt_add[3]~11_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_add[3]~12 ;
//wire	\eth_udp_inst|ip_send_inst|cnt_add [4];
wire	\eth_udp_inst|ip_send_inst|cnt_add[4]~13_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_add[4]~15_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout ;
wire	[2:0] \eth_udp_inst|ip_send_inst|cnt_send_bit ;
//wire	\eth_udp_inst|ip_send_inst|cnt_send_bit [0];
//wire	\eth_udp_inst|ip_send_inst|cnt_send_bit [1];
//wire	\eth_udp_inst|ip_send_inst|cnt_send_bit [2];
wire	\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_send_bit~2_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_send_bit~4_combout ;
wire	\eth_udp_inst|ip_send_inst|cnt_send_bit~5_combout ;
wire	\eth_udp_inst|ip_send_inst|crc_clr~q ;
wire	\eth_udp_inst|ip_send_inst|crc_en~q ;
wire	[15:0] \eth_udp_inst|ip_send_inst|data_cnt ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [0];
wire	\eth_udp_inst|ip_send_inst|data_cnt[0]~16_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[0]~17 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [10];
wire	\eth_udp_inst|ip_send_inst|data_cnt[10]~36_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[10]~37 ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [11];
wire	\eth_udp_inst|ip_send_inst|data_cnt[11]~42_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[11]~43 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [12];
wire	\eth_udp_inst|ip_send_inst|data_cnt[12]~44_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[12]~45 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [13];
wire	\eth_udp_inst|ip_send_inst|data_cnt[13]~46_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[13]~47 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [14];
wire	\eth_udp_inst|ip_send_inst|data_cnt[14]~48_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[14]~49 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [15];
wire	\eth_udp_inst|ip_send_inst|data_cnt[15]~50_combout ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [1];
wire	\eth_udp_inst|ip_send_inst|data_cnt[1]~18_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[1]~19 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [2];
wire	\eth_udp_inst|ip_send_inst|data_cnt[2]~20_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[2]~21 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [3];
wire	\eth_udp_inst|ip_send_inst|data_cnt[3]~22_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[3]~23 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [4];
wire	\eth_udp_inst|ip_send_inst|data_cnt[4]~24_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[4]~25 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [5];
wire	\eth_udp_inst|ip_send_inst|data_cnt[5]~26_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[5]~27 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [6];
wire	\eth_udp_inst|ip_send_inst|data_cnt[6]~28_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[6]~29 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [7];
wire	\eth_udp_inst|ip_send_inst|data_cnt[7]~30_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[7]~31 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [8];
wire	\eth_udp_inst|ip_send_inst|data_cnt[8]~32_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[8]~33 ;
//wire	\eth_udp_inst|ip_send_inst|data_cnt [9];
wire	\eth_udp_inst|ip_send_inst|data_cnt[9]~34_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[9]~35 ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[9]~38_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[9]~39_combout ;
wire	\eth_udp_inst|ip_send_inst|data_cnt[9]~40_combout ;
wire	[15:0] \eth_udp_inst|ip_send_inst|data_len ;
//wire	\eth_udp_inst|ip_send_inst|data_len [0];
//wire	\eth_udp_inst|ip_send_inst|data_len [10];
wire	\eth_udp_inst|ip_send_inst|data_len[10]~0_combout ;
//wire	\eth_udp_inst|ip_send_inst|data_len [11];
//wire	\eth_udp_inst|ip_send_inst|data_len [12];
//wire	\eth_udp_inst|ip_send_inst|data_len [13];
//wire	\eth_udp_inst|ip_send_inst|data_len [14];
//wire	\eth_udp_inst|ip_send_inst|data_len [15];
//wire	\eth_udp_inst|ip_send_inst|data_len [1];
//wire	\eth_udp_inst|ip_send_inst|data_len [2];
//wire	\eth_udp_inst|ip_send_inst|data_len [3];
//wire	\eth_udp_inst|ip_send_inst|data_len [4];
//wire	\eth_udp_inst|ip_send_inst|data_len [5];
//wire	\eth_udp_inst|ip_send_inst|data_len [6];
//wire	\eth_udp_inst|ip_send_inst|data_len [7];
//wire	\eth_udp_inst|ip_send_inst|data_len [8];
//wire	\eth_udp_inst|ip_send_inst|data_len [9];
wire	[3:0] \eth_udp_inst|ip_send_inst|eth_tx_data ;
//wire	\eth_udp_inst|ip_send_inst|eth_tx_data [0];
//wire	\eth_udp_inst|ip_send_inst|eth_tx_data [1];
//wire	\eth_udp_inst|ip_send_inst|eth_tx_data [2];
//wire	\eth_udp_inst|ip_send_inst|eth_tx_data [3];
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~0_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~10_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~11_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~12_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~13_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~14_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~15_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~16_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~17_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~18_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~19_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~1_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~20_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~21_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~22_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~23_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~24_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~25_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~26_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~27_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~28_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~29_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~2_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~30_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~31_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~32_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~33_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~34_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~35_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~36_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~37_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~38_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~39_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~3_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~40_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~41_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~42_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~43_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~44_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~45_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~46_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~47_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~48_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~49_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~4_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~50_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~51_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~52_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~53_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~54_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~55_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~56_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~57_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~58_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~59_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~5_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~60_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~61_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~62_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~63_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~64_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~65_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~66_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~67_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~68_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~69_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~6_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~70_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~71_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~72_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~73_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~74_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~75_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~76_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~77_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~78_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~79_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~7_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~80_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~81_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~82_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~83_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~84_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~85_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~86_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~87_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~88_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~89_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~8_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~90_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~91_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_data~9_combout ;
wire	\eth_udp_inst|ip_send_inst|eth_tx_en~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~18_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~53_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~21_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~22 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~23_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~24 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~25_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~26 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~27_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~28 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~29_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~30 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~31_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~32 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~33_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~34 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~35_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~36 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~37_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~38 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~39_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~40 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~41_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~42 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~43_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~44 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~45_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~46 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~47_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~48 ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~58_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][0]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][10]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][11]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][12]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][13]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][14]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][15]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][1]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][2]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][3]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][4]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][5]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][6]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][7]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head[2][9]~q ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~15_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~17_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~19_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~20_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~49_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~50_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~51_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~52_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~54_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~55_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~56_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~57_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~60_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~61_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~62_combout ;
wire	\eth_udp_inst|ip_send_inst|ip_udp_head~63_combout ;
wire	\eth_udp_inst|ip_send_inst|packet_head[7][7]~feeder_combout ;
wire	\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ;
wire	\eth_udp_inst|ip_send_inst|read_data_req~0_combout ;
wire	\eth_udp_inst|ip_send_inst|read_data_req~q ;
wire	\eth_udp_inst|ip_send_inst|send_en_r~q ;
wire	\eth_udp_inst|ip_send_inst|send_end~q ;
wire	\eth_udp_inst|ip_send_inst|state.CHECK_SUM~0_combout ;
wire	\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ;
wire	\eth_udp_inst|ip_send_inst|state.CRC~q ;
wire	\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ;
wire	\eth_udp_inst|ip_send_inst|state.IDLE~0_combout ;
wire	\eth_udp_inst|ip_send_inst|state.IDLE~q ;
wire	\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ;
wire	\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ;
wire	\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ;
wire	\eth_udp_inst|ip_send_inst|sw_en~0_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~1_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~2_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~3_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~4_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~5_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~6_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~7_combout ;
wire	\eth_udp_inst|ip_send_inst|sw_en~q ;
wire	\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ;
wire	\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y16_SIG ;
wire	\led_r~0_combout ;
wire	\led_r~q ;
wire	[1:0] \mii_to_rmii_inst|eth_tx_data ;
//wire	\mii_to_rmii_inst|eth_tx_data [0];
wire	\mii_to_rmii_inst|eth_tx_data[0]~feeder_combout ;
//wire	\mii_to_rmii_inst|eth_tx_data [1];
wire	\mii_to_rmii_inst|eth_tx_data[1]~feeder_combout ;
wire	[1:0] \mii_to_rmii_inst|eth_tx_data_reg ;
//wire	\mii_to_rmii_inst|eth_tx_data_reg [0];
//wire	\mii_to_rmii_inst|eth_tx_data_reg [1];
wire	\mii_to_rmii_inst|eth_tx_data_reg~0_combout ;
wire	\mii_to_rmii_inst|eth_tx_data_reg~1_combout ;
wire	\mii_to_rmii_inst|eth_tx_dv~feeder_combout ;
wire	\mii_to_rmii_inst|eth_tx_dv~q ;
wire	\mii_to_rmii_inst|rd_flag~0_combout ;
wire	\mii_to_rmii_inst|rd_flag~q ;
wire	[3:0] \mii_to_rmii_inst|tx_data_reg ;
//wire	\mii_to_rmii_inst|tx_data_reg [0];
wire	\mii_to_rmii_inst|tx_data_reg[0]~feeder_combout ;
//wire	\mii_to_rmii_inst|tx_data_reg [1];
//wire	\mii_to_rmii_inst|tx_data_reg [2];
wire	\mii_to_rmii_inst|tx_data_reg[2]~feeder_combout ;
//wire	\mii_to_rmii_inst|tx_data_reg [3];
wire	\mii_to_rmii_inst|tx_data_reg[3]~feeder_combout ;
wire	\mii_to_rmii_inst|tx_dv_reg~feeder_combout ;
wire	\mii_to_rmii_inst|tx_dv_reg~q ;
wire	[5:0] reset_init;
//wire	reset_init[0];
wire	\reset_init[0]~1_combout ;
//wire	reset_init[1];
//wire	reset_init[2];
//wire	reset_init[3];
//wire	reset_init[4];
//wire	reset_init[5];
wire	\reset_init[5]~0_combout ;
wire	\reset_init[5]~clkctrl_outclk ;
wire	\reset_init[5]~clkctrl_outclk__AsyncReset_X1_Y1_INV ;
wire	\rst_n~input_o ;
wire	[24:0] timer;
//wire	timer[0];
wire	\timer[0]~25_combout ;
wire	\timer[0]~26 ;
//wire	timer[10];
wire	\timer[10]~45_combout ;
wire	\timer[10]~46 ;
//wire	timer[11];
wire	\timer[11]~47_combout ;
wire	\timer[11]~48 ;
//wire	timer[12];
wire	\timer[12]~49_combout ;
wire	\timer[12]~50 ;
//wire	timer[13];
wire	\timer[13]~51_combout ;
wire	\timer[13]~52 ;
//wire	timer[14];
wire	\timer[14]~53_combout ;
wire	\timer[14]~54 ;
//wire	timer[15];
wire	\timer[15]~55_combout ;
wire	\timer[15]~56 ;
//wire	timer[16];
wire	\timer[16]~57_combout ;
wire	\timer[16]~58 ;
//wire	timer[17];
wire	\timer[17]~59_combout ;
wire	\timer[17]~60 ;
//wire	timer[18];
wire	\timer[18]~61_combout ;
wire	\timer[18]~62 ;
//wire	timer[19];
wire	\timer[19]~63_combout ;
wire	\timer[19]~64 ;
//wire	timer[1];
wire	\timer[1]~27_combout ;
wire	\timer[1]~28 ;
//wire	timer[20];
wire	\timer[20]~65_combout ;
wire	\timer[20]~66 ;
//wire	timer[21];
wire	\timer[21]~67_combout ;
wire	\timer[21]~68 ;
//wire	timer[22];
wire	\timer[22]~69_combout ;
wire	\timer[22]~70 ;
//wire	timer[23];
wire	\timer[23]~71_combout ;
wire	\timer[23]~72 ;
//wire	timer[24];
wire	\timer[24]~73_combout ;
//wire	timer[2];
wire	\timer[2]~29_combout ;
wire	\timer[2]~30 ;
//wire	timer[3];
wire	\timer[3]~31_combout ;
wire	\timer[3]~32 ;
//wire	timer[4];
wire	\timer[4]~33_combout ;
wire	\timer[4]~34 ;
//wire	timer[5];
wire	\timer[5]~35_combout ;
wire	\timer[5]~36 ;
//wire	timer[6];
wire	\timer[6]~37_combout ;
wire	\timer[6]~38 ;
//wire	timer[7];
wire	\timer[7]~39_combout ;
wire	\timer[7]~40 ;
//wire	timer[8];
wire	\timer[8]~41_combout ;
wire	\timer[8]~42 ;
//wire	timer[9];
wire	\timer[9]~43_combout ;
wire	\timer[9]~44 ;
wire	unknown;
wire	\~QIC_CREATED_GND~I_combout ;

wire vcc;
wire gnd;
assign vcc = 1'b1;
assign gnd = 1'b0;

alta_slice \Add0~8 (
	.A(vcc),
	.B(reset_init[5]),
	.C(vcc),
	.D(vcc),
	.Cin(\Add0~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Add0~8_combout ),
	.Cout(),
	.Q());
defparam \Add0~8 .coord_x = 47;
defparam \Add0~8 .coord_y = 15;
defparam \Add0~8 .coord_z = 9;
defparam \Add0~8 .mask = 16'hC3C3;
defparam \Add0~8 .modeMux = 1'b1;
defparam \Add0~8 .FeedbackMux = 1'b0;
defparam \Add0~8 .ShiftMux = 1'b0;
defparam \Add0~8 .BypassEn = 1'b0;
defparam \Add0~8 .CarryEnb = 1'b1;

alta_slice \Equal0~0 (
	.A(timer[1]),
	.B(timer[0]),
	.C(timer[3]),
	.D(timer[2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~0_combout ),
	.Cout(),
	.Q());
defparam \Equal0~0 .coord_x = 2;
defparam \Equal0~0 .coord_y = 12;
defparam \Equal0~0 .coord_z = 0;
defparam \Equal0~0 .mask = 16'h0001;
defparam \Equal0~0 .modeMux = 1'b0;
defparam \Equal0~0 .FeedbackMux = 1'b0;
defparam \Equal0~0 .ShiftMux = 1'b0;
defparam \Equal0~0 .BypassEn = 1'b0;
defparam \Equal0~0 .CarryEnb = 1'b1;

alta_slice \Equal0~1 (
	.A(timer[7]),
	.B(timer[5]),
	.C(timer[4]),
	.D(timer[6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~1_combout ),
	.Cout(),
	.Q());
defparam \Equal0~1 .coord_x = 2;
defparam \Equal0~1 .coord_y = 12;
defparam \Equal0~1 .coord_z = 1;
defparam \Equal0~1 .mask = 16'h0001;
defparam \Equal0~1 .modeMux = 1'b0;
defparam \Equal0~1 .FeedbackMux = 1'b0;
defparam \Equal0~1 .ShiftMux = 1'b0;
defparam \Equal0~1 .BypassEn = 1'b0;
defparam \Equal0~1 .CarryEnb = 1'b1;

alta_slice \Equal0~2 (
	.A(timer[11]),
	.B(timer[8]),
	.C(timer[10]),
	.D(timer[9]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~2_combout ),
	.Cout(),
	.Q());
defparam \Equal0~2 .coord_x = 2;
defparam \Equal0~2 .coord_y = 12;
defparam \Equal0~2 .coord_z = 2;
defparam \Equal0~2 .mask = 16'h0001;
defparam \Equal0~2 .modeMux = 1'b0;
defparam \Equal0~2 .FeedbackMux = 1'b0;
defparam \Equal0~2 .ShiftMux = 1'b0;
defparam \Equal0~2 .BypassEn = 1'b0;
defparam \Equal0~2 .CarryEnb = 1'b1;

alta_slice \Equal0~3 (
	.A(timer[12]),
	.B(timer[14]),
	.C(timer[13]),
	.D(timer[15]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~3_combout ),
	.Cout(),
	.Q());
defparam \Equal0~3 .coord_x = 2;
defparam \Equal0~3 .coord_y = 11;
defparam \Equal0~3 .coord_z = 13;
defparam \Equal0~3 .mask = 16'h0001;
defparam \Equal0~3 .modeMux = 1'b0;
defparam \Equal0~3 .FeedbackMux = 1'b0;
defparam \Equal0~3 .ShiftMux = 1'b0;
defparam \Equal0~3 .BypassEn = 1'b0;
defparam \Equal0~3 .CarryEnb = 1'b1;

alta_slice \Equal0~4 (
	.A(\Equal0~0_combout ),
	.B(\Equal0~2_combout ),
	.C(\Equal0~1_combout ),
	.D(\Equal0~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~4_combout ),
	.Cout(),
	.Q());
defparam \Equal0~4 .coord_x = 2;
defparam \Equal0~4 .coord_y = 12;
defparam \Equal0~4 .coord_z = 3;
defparam \Equal0~4 .mask = 16'h8000;
defparam \Equal0~4 .modeMux = 1'b0;
defparam \Equal0~4 .FeedbackMux = 1'b0;
defparam \Equal0~4 .ShiftMux = 1'b0;
defparam \Equal0~4 .BypassEn = 1'b0;
defparam \Equal0~4 .CarryEnb = 1'b1;

alta_slice \Equal0~5 (
	.A(timer[17]),
	.B(timer[16]),
	.C(timer[19]),
	.D(timer[18]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~5_combout ),
	.Cout(),
	.Q());
defparam \Equal0~5 .coord_x = 2;
defparam \Equal0~5 .coord_y = 11;
defparam \Equal0~5 .coord_z = 14;
defparam \Equal0~5 .mask = 16'h0001;
defparam \Equal0~5 .modeMux = 1'b0;
defparam \Equal0~5 .FeedbackMux = 1'b0;
defparam \Equal0~5 .ShiftMux = 1'b0;
defparam \Equal0~5 .BypassEn = 1'b0;
defparam \Equal0~5 .CarryEnb = 1'b1;

alta_slice \Equal0~6 (
	.A(timer[23]),
	.B(timer[20]),
	.C(timer[22]),
	.D(timer[21]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~6_combout ),
	.Cout(),
	.Q());
defparam \Equal0~6 .coord_x = 2;
defparam \Equal0~6 .coord_y = 11;
defparam \Equal0~6 .coord_z = 15;
defparam \Equal0~6 .mask = 16'h0001;
defparam \Equal0~6 .modeMux = 1'b0;
defparam \Equal0~6 .FeedbackMux = 1'b0;
defparam \Equal0~6 .ShiftMux = 1'b0;
defparam \Equal0~6 .BypassEn = 1'b0;
defparam \Equal0~6 .CarryEnb = 1'b1;

alta_slice \Equal0~7 (
	.A(vcc),
	.B(vcc),
	.C(\Equal0~6_combout ),
	.D(timer[24]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Equal0~7_combout ),
	.Cout(),
	.Q());
defparam \Equal0~7 .coord_x = 1;
defparam \Equal0~7 .coord_y = 11;
defparam \Equal0~7 .coord_z = 8;
defparam \Equal0~7 .mask = 16'h00F0;
defparam \Equal0~7 .modeMux = 1'b0;
defparam \Equal0~7 .FeedbackMux = 1'b0;
defparam \Equal0~7 .ShiftMux = 1'b0;
defparam \Equal0~7 .BypassEn = 1'b0;
defparam \Equal0~7 .CarryEnb = 1'b1;

alta_slice \alt_pll_inst|altpll_component|auto_generated|locked (
	.A(\alt_pll_inst|altpll_component|auto_generated|pll_lock_sync~q ),
	.B(vcc),
	.C(vcc),
	.D(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.Cout(),
	.Q());
defparam \alt_pll_inst|altpll_component|auto_generated|locked .coord_x = 1;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .coord_y = 12;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .coord_z = 11;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .mask = 16'h55FF;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .modeMux = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .FeedbackMux = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .ShiftMux = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .BypassEn = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|locked .CarryEnb = 1'b1;

alta_io_gclk \alt_pll_inst|altpll_component|auto_generated|locked~clkctrl (
	.inclk(\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.outclk(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ));
defparam \alt_pll_inst|altpll_component|auto_generated|locked~clkctrl .coord_x = 0;
defparam \alt_pll_inst|altpll_component|auto_generated|locked~clkctrl .coord_y = 12;
defparam \alt_pll_inst|altpll_component|auto_generated|locked~clkctrl .coord_z = 2;

alta_pllve \alt_pll_inst|altpll_component|auto_generated|pll1 (
	.clkin(\clk~input_o ),
	.clkfb(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_fbout ),
	.pfden(vcc),
	.resetn(\reset_init[5]~clkctrl_outclk ),
	.phasecounterselect({gnd, gnd, gnd}),
	.phaseupdown(gnd),
	.phasestep(gnd),
	.scanclk(gnd),
	.scanclkena(vcc),
	.scandata(gnd),
	.configupdate(gnd),
	.scandataout(),
	.scandone(),
	.phasedone(),
	.clkout0(\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [0]),
	.clkout1(\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [1]),
	.clkout2(\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [2]),
	.clkout3(\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [3]),
	.clkout4(\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [4]),
	.clkfbout(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_fbout ),
	.lock(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked ));
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .coord_x = 0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .coord_y = 1;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .coord_z = 0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKIN_HIGH = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKIN_LOW = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKIN_TRIM = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKIN_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKFB_HIGH = 8'b00010001;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKFB_LOW = 8'b00010010;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKFB_TRIM = 1'b1;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKFB_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKDIV0_EN = 1'b1;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKDIV1_EN = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKDIV2_EN = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKDIV3_EN = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKDIV4_EN = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT0_HIGH = 8'b00010001;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT0_LOW = 8'b00010010;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT0_TRIM = 1'b1;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT0_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_HIGH = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_LOW = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_TRIM = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_HIGH = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_LOW = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_TRIM = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_HIGH = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_LOW = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_TRIM = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_HIGH = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_LOW = 8'b11111111;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_TRIM = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_BYPASS = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT0_DEL = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_DEL = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_DEL = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_DEL = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_DEL = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT0_PHASE = 3'b000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_PHASE = 3'b000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_PHASE = 3'b000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_PHASE = 3'b000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_PHASE = 3'b000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKFB_DEL = 8'b00000000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKFB_PHASE = 3'b000;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .FEEDBACK_MODE = 3'b100;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .FBDELAY_VAL = 3'b100;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .PLLOUTP_EN = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .PLLOUTN_EN = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT1_CASCADE = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT2_CASCADE = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT3_CASCADE = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CLKOUT4_CASCADE = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .VCO_POST_DIV = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .REG_CTRL = 2'b10;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .CP = 3'b100;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .RREF = 2'b01;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .RVI = 2'b01;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .IVCO = 3'b010;
defparam \alt_pll_inst|altpll_component|auto_generated|pll1 .PLL_EN_FLAG = 1'b1;

alta_slice \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\alt_pll_inst|altpll_component|auto_generated|pll_lock_sync~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked_X1_Y1_SIG_VCC ),
	.AsyncReset(\reset_init[5]~clkctrl_outclk__AsyncReset_X1_Y1_INV ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\alt_pll_inst|altpll_component|auto_generated|pll_lock_sync~feeder_combout ),
	.Cout(),
	.Q(\alt_pll_inst|altpll_component|auto_generated|pll_lock_sync~q ));
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .coord_x = 1;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .coord_y = 12;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .coord_z = 15;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .mask = 16'hFFFF;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .modeMux = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .FeedbackMux = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .ShiftMux = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .BypassEn = 1'b0;
defparam \alt_pll_inst|altpll_component|auto_generated|pll_lock_sync .CarryEnb = 1'b1;

alta_io_gclk \alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl (
	.inclk(\alt_pll_inst|altpll_component|auto_generated|pll1_CLK_bus [0]),
	.outclk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ));
defparam \alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl .coord_x = 0;
defparam \alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl .coord_y = 12;
defparam \alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl .coord_z = 3;

alta_jtag altera_internal_jtag(
	.tdouser(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());
defparam altera_internal_jtag.coord_x = 1;
defparam altera_internal_jtag.coord_y = 18;
defparam altera_internal_jtag.coord_z = 0;

alta_io_gclk \altera_internal_jtag~TCKUTAPclkctrl (
	.inclk(\altera_internal_jtag~TCKUTAP ),
	.outclk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ));
defparam \altera_internal_jtag~TCKUTAPclkctrl .coord_x = 0;
defparam \altera_internal_jtag~TCKUTAPclkctrl .coord_y = 12;
defparam \altera_internal_jtag~TCKUTAPclkctrl .coord_z = 1;

alta_asyncctrl asyncreset_ctrl_X10_Y9_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ));
defparam asyncreset_ctrl_X10_Y9_N0.coord_x = 16;
defparam asyncreset_ctrl_X10_Y9_N0.coord_y = 13;
defparam asyncreset_ctrl_X10_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X10_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X11_Y14_N0(
	.Din(),
	.Dout(AsyncReset_X11_Y14_GND));
defparam asyncreset_ctrl_X11_Y14_N0.coord_x = 9;
defparam asyncreset_ctrl_X11_Y14_N0.coord_y = 14;
defparam asyncreset_ctrl_X11_Y14_N0.coord_z = 0;
defparam asyncreset_ctrl_X11_Y14_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X11_Y14_N1(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X11_Y14_SIG ));
defparam asyncreset_ctrl_X11_Y14_N1.coord_x = 9;
defparam asyncreset_ctrl_X11_Y14_N1.coord_y = 14;
defparam asyncreset_ctrl_X11_Y14_N1.coord_z = 1;
defparam asyncreset_ctrl_X11_Y14_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X11_Y16_N0(
	.Din(),
	.Dout(AsyncReset_X11_Y16_GND));
defparam asyncreset_ctrl_X11_Y16_N0.coord_x = 16;
defparam asyncreset_ctrl_X11_Y16_N0.coord_y = 15;
defparam asyncreset_ctrl_X11_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X11_Y16_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X11_Y9_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ));
defparam asyncreset_ctrl_X11_Y9_N0.coord_x = 16;
defparam asyncreset_ctrl_X11_Y9_N0.coord_y = 12;
defparam asyncreset_ctrl_X11_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X11_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X12_Y14_N0(
	.Din(),
	.Dout(AsyncReset_X12_Y14_GND));
defparam asyncreset_ctrl_X12_Y14_N0.coord_x = 10;
defparam asyncreset_ctrl_X12_Y14_N0.coord_y = 14;
defparam asyncreset_ctrl_X12_Y14_N0.coord_z = 0;
defparam asyncreset_ctrl_X12_Y14_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X12_Y14_N1(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y14_SIG ));
defparam asyncreset_ctrl_X12_Y14_N1.coord_x = 10;
defparam asyncreset_ctrl_X12_Y14_N1.coord_y = 14;
defparam asyncreset_ctrl_X12_Y14_N1.coord_z = 1;
defparam asyncreset_ctrl_X12_Y14_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X12_Y16_N0(
	.Din(),
	.Dout(AsyncReset_X12_Y16_GND));
defparam asyncreset_ctrl_X12_Y16_N0.coord_x = 17;
defparam asyncreset_ctrl_X12_Y16_N0.coord_y = 15;
defparam asyncreset_ctrl_X12_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X12_Y16_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X12_Y18_N0(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y18_SIG ));
defparam asyncreset_ctrl_X12_Y18_N0.coord_x = 11;
defparam asyncreset_ctrl_X12_Y18_N0.coord_y = 14;
defparam asyncreset_ctrl_X12_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X12_Y18_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X12_Y18_N1(
	.Din(),
	.Dout(AsyncReset_X12_Y18_GND));
defparam asyncreset_ctrl_X12_Y18_N1.coord_x = 11;
defparam asyncreset_ctrl_X12_Y18_N1.coord_y = 14;
defparam asyncreset_ctrl_X12_Y18_N1.coord_z = 1;
defparam asyncreset_ctrl_X12_Y18_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X12_Y9_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y9_SIG ));
defparam asyncreset_ctrl_X12_Y9_N0.coord_x = 15;
defparam asyncreset_ctrl_X12_Y9_N0.coord_y = 11;
defparam asyncreset_ctrl_X12_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X12_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X13_Y10_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y10_SIG ));
defparam asyncreset_ctrl_X13_Y10_N0.coord_x = 17;
defparam asyncreset_ctrl_X13_Y10_N0.coord_y = 12;
defparam asyncreset_ctrl_X13_Y10_N0.coord_z = 0;
defparam asyncreset_ctrl_X13_Y10_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X13_Y16_N0(
	.Din(),
	.Dout(AsyncReset_X13_Y16_GND));
defparam asyncreset_ctrl_X13_Y16_N0.coord_x = 17;
defparam asyncreset_ctrl_X13_Y16_N0.coord_y = 14;
defparam asyncreset_ctrl_X13_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X13_Y16_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X13_Y18_N0(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X13_Y18_SIG ));
defparam asyncreset_ctrl_X13_Y18_N0.coord_x = 10;
defparam asyncreset_ctrl_X13_Y18_N0.coord_y = 12;
defparam asyncreset_ctrl_X13_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X13_Y18_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X13_Y18_N1(
	.Din(),
	.Dout(AsyncReset_X13_Y18_GND));
defparam asyncreset_ctrl_X13_Y18_N1.coord_x = 10;
defparam asyncreset_ctrl_X13_Y18_N1.coord_y = 12;
defparam asyncreset_ctrl_X13_Y18_N1.coord_z = 1;
defparam asyncreset_ctrl_X13_Y18_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X13_Y7_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y7_SIG ));
defparam asyncreset_ctrl_X13_Y7_N0.coord_x = 17;
defparam asyncreset_ctrl_X13_Y7_N0.coord_y = 13;
defparam asyncreset_ctrl_X13_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X13_Y7_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X13_Y9_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ));
defparam asyncreset_ctrl_X13_Y9_N0.coord_x = 16;
defparam asyncreset_ctrl_X13_Y9_N0.coord_y = 11;
defparam asyncreset_ctrl_X13_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X13_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X14_Y10_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ));
defparam asyncreset_ctrl_X14_Y10_N0.coord_x = 16;
defparam asyncreset_ctrl_X14_Y10_N0.coord_y = 9;
defparam asyncreset_ctrl_X14_Y10_N0.coord_z = 0;
defparam asyncreset_ctrl_X14_Y10_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X14_Y11_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y11_SIG ));
defparam asyncreset_ctrl_X14_Y11_N0.coord_x = 15;
defparam asyncreset_ctrl_X14_Y11_N0.coord_y = 10;
defparam asyncreset_ctrl_X14_Y11_N0.coord_z = 0;
defparam asyncreset_ctrl_X14_Y11_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X14_Y14_N0(
	.Din(),
	.Dout(AsyncReset_X14_Y14_GND));
defparam asyncreset_ctrl_X14_Y14_N0.coord_x = 14;
defparam asyncreset_ctrl_X14_Y14_N0.coord_y = 15;
defparam asyncreset_ctrl_X14_Y14_N0.coord_z = 0;
defparam asyncreset_ctrl_X14_Y14_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X14_Y16_N0(
	.Din(),
	.Dout(AsyncReset_X14_Y16_GND));
defparam asyncreset_ctrl_X14_Y16_N0.coord_x = 13;
defparam asyncreset_ctrl_X14_Y16_N0.coord_y = 14;
defparam asyncreset_ctrl_X14_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X14_Y16_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X14_Y18_N0(
	.Din(),
	.Dout(AsyncReset_X14_Y18_GND));
defparam asyncreset_ctrl_X14_Y18_N0.coord_x = 13;
defparam asyncreset_ctrl_X14_Y18_N0.coord_y = 12;
defparam asyncreset_ctrl_X14_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X14_Y18_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X14_Y19_N0(
	.Din(),
	.Dout(AsyncReset_X14_Y19_GND));
defparam asyncreset_ctrl_X14_Y19_N0.coord_x = 8;
defparam asyncreset_ctrl_X14_Y19_N0.coord_y = 9;
defparam asyncreset_ctrl_X14_Y19_N0.coord_z = 0;
defparam asyncreset_ctrl_X14_Y19_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X14_Y20_N0(
	.Din(),
	.Dout(AsyncReset_X14_Y20_GND));
defparam asyncreset_ctrl_X14_Y20_N0.coord_x = 8;
defparam asyncreset_ctrl_X14_Y20_N0.coord_y = 10;
defparam asyncreset_ctrl_X14_Y20_N0.coord_z = 0;
defparam asyncreset_ctrl_X14_Y20_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X14_Y8_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ));
defparam asyncreset_ctrl_X14_Y8_N0.coord_x = 16;
defparam asyncreset_ctrl_X14_Y8_N0.coord_y = 10;
defparam asyncreset_ctrl_X14_Y8_N0.coord_z = 0;
defparam asyncreset_ctrl_X14_Y8_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X14_Y9_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y9_SIG ));
defparam asyncreset_ctrl_X14_Y9_N0.coord_x = 17;
defparam asyncreset_ctrl_X14_Y9_N0.coord_y = 11;
defparam asyncreset_ctrl_X14_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X14_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X16_Y10_N0(
	.Din(),
	.Dout(AsyncReset_X16_Y10_GND));
defparam asyncreset_ctrl_X16_Y10_N0.coord_x = 19;
defparam asyncreset_ctrl_X16_Y10_N0.coord_y = 9;
defparam asyncreset_ctrl_X16_Y10_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y10_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X16_Y11_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y11_SIG ));
defparam asyncreset_ctrl_X16_Y11_N0.coord_x = 20;
defparam asyncreset_ctrl_X16_Y11_N0.coord_y = 5;
defparam asyncreset_ctrl_X16_Y11_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y11_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X16_Y12_N0(
	.Din(),
	.Dout(AsyncReset_X16_Y12_GND));
defparam asyncreset_ctrl_X16_Y12_N0.coord_x = 19;
defparam asyncreset_ctrl_X16_Y12_N0.coord_y = 11;
defparam asyncreset_ctrl_X16_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y12_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X16_Y14_N0(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ));
defparam asyncreset_ctrl_X16_Y14_N0.coord_x = 13;
defparam asyncreset_ctrl_X16_Y14_N0.coord_y = 15;
defparam asyncreset_ctrl_X16_Y14_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y14_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X16_Y16_N0(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ));
defparam asyncreset_ctrl_X16_Y16_N0.coord_x = 15;
defparam asyncreset_ctrl_X16_Y16_N0.coord_y = 15;
defparam asyncreset_ctrl_X16_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y16_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X16_Y16_N1(
	.Din(),
	.Dout(AsyncReset_X16_Y16_GND));
defparam asyncreset_ctrl_X16_Y16_N1.coord_x = 15;
defparam asyncreset_ctrl_X16_Y16_N1.coord_y = 15;
defparam asyncreset_ctrl_X16_Y16_N1.coord_z = 1;
defparam asyncreset_ctrl_X16_Y16_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X16_Y17_N0(
	.Din(),
	.Dout(AsyncReset_X16_Y17_GND));
defparam asyncreset_ctrl_X16_Y17_N0.coord_x = 17;
defparam asyncreset_ctrl_X16_Y17_N0.coord_y = 16;
defparam asyncreset_ctrl_X16_Y17_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y17_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X16_Y18_N0(
	.Din(),
	.Dout(AsyncReset_X16_Y18_GND));
defparam asyncreset_ctrl_X16_Y18_N0.coord_x = 14;
defparam asyncreset_ctrl_X16_Y18_N0.coord_y = 14;
defparam asyncreset_ctrl_X16_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y18_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X16_Y19_N0(
	.Din(),
	.Dout(AsyncReset_X16_Y19_GND));
defparam asyncreset_ctrl_X16_Y19_N0.coord_x = 14;
defparam asyncreset_ctrl_X16_Y19_N0.coord_y = 12;
defparam asyncreset_ctrl_X16_Y19_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y19_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X16_Y8_N0(
	.Din(),
	.Dout(AsyncReset_X16_Y8_GND));
defparam asyncreset_ctrl_X16_Y8_N0.coord_x = 17;
defparam asyncreset_ctrl_X16_Y8_N0.coord_y = 10;
defparam asyncreset_ctrl_X16_Y8_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y8_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X16_Y8_N1(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y8_SIG ));
defparam asyncreset_ctrl_X16_Y8_N1.coord_x = 17;
defparam asyncreset_ctrl_X16_Y8_N1.coord_y = 10;
defparam asyncreset_ctrl_X16_Y8_N1.coord_z = 1;
defparam asyncreset_ctrl_X16_Y8_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X16_Y9_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ));
defparam asyncreset_ctrl_X16_Y9_N0.coord_x = 17;
defparam asyncreset_ctrl_X16_Y9_N0.coord_y = 9;
defparam asyncreset_ctrl_X16_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X16_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X17_Y10_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y10_SIG ));
defparam asyncreset_ctrl_X17_Y10_N0.coord_x = 24;
defparam asyncreset_ctrl_X17_Y10_N0.coord_y = 6;
defparam asyncreset_ctrl_X17_Y10_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y10_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X17_Y11_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y11_SIG ));
defparam asyncreset_ctrl_X17_Y11_N0.coord_x = 24;
defparam asyncreset_ctrl_X17_Y11_N0.coord_y = 5;
defparam asyncreset_ctrl_X17_Y11_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y11_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X17_Y14_N0(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ));
defparam asyncreset_ctrl_X17_Y14_N0.coord_x = 12;
defparam asyncreset_ctrl_X17_Y14_N0.coord_y = 15;
defparam asyncreset_ctrl_X17_Y14_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y14_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X17_Y15_N0(
	.Din(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.Dout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X17_Y15_SIG ));
defparam asyncreset_ctrl_X17_Y15_N0.coord_x = 5;
defparam asyncreset_ctrl_X17_Y15_N0.coord_y = 15;
defparam asyncreset_ctrl_X17_Y15_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y15_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X17_Y15_N1(
	.Din(),
	.Dout(AsyncReset_X17_Y15_GND));
defparam asyncreset_ctrl_X17_Y15_N1.coord_x = 5;
defparam asyncreset_ctrl_X17_Y15_N1.coord_y = 15;
defparam asyncreset_ctrl_X17_Y15_N1.coord_z = 1;
defparam asyncreset_ctrl_X17_Y15_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X17_Y16_N0(
	.Din(),
	.Dout(AsyncReset_X17_Y16_GND));
defparam asyncreset_ctrl_X17_Y16_N0.coord_x = 7;
defparam asyncreset_ctrl_X17_Y16_N0.coord_y = 17;
defparam asyncreset_ctrl_X17_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y16_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X17_Y17_N0(
	.Din(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.Dout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X17_Y17_SIG ));
defparam asyncreset_ctrl_X17_Y17_N0.coord_x = 6;
defparam asyncreset_ctrl_X17_Y17_N0.coord_y = 16;
defparam asyncreset_ctrl_X17_Y17_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y17_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X17_Y18_N0(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y18_SIG ));
defparam asyncreset_ctrl_X17_Y18_N0.coord_x = 15;
defparam asyncreset_ctrl_X17_Y18_N0.coord_y = 14;
defparam asyncreset_ctrl_X17_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y18_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X17_Y18_N1(
	.Din(),
	.Dout(AsyncReset_X17_Y18_GND));
defparam asyncreset_ctrl_X17_Y18_N1.coord_x = 15;
defparam asyncreset_ctrl_X17_Y18_N1.coord_y = 14;
defparam asyncreset_ctrl_X17_Y18_N1.coord_z = 1;
defparam asyncreset_ctrl_X17_Y18_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X17_Y19_N0(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y19_SIG ));
defparam asyncreset_ctrl_X17_Y19_N0.coord_x = 15;
defparam asyncreset_ctrl_X17_Y19_N0.coord_y = 12;
defparam asyncreset_ctrl_X17_Y19_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y19_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X17_Y19_N1(
	.Din(),
	.Dout(AsyncReset_X17_Y19_GND));
defparam asyncreset_ctrl_X17_Y19_N1.coord_x = 15;
defparam asyncreset_ctrl_X17_Y19_N1.coord_y = 12;
defparam asyncreset_ctrl_X17_Y19_N1.coord_z = 1;
defparam asyncreset_ctrl_X17_Y19_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X17_Y20_N0(
	.Din(),
	.Dout(AsyncReset_X17_Y20_GND));
defparam asyncreset_ctrl_X17_Y20_N0.coord_x = 14;
defparam asyncreset_ctrl_X17_Y20_N0.coord_y = 16;
defparam asyncreset_ctrl_X17_Y20_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y20_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X17_Y9_N0(
	.Din(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.Dout(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ));
defparam asyncreset_ctrl_X17_Y9_N0.coord_x = 15;
defparam asyncreset_ctrl_X17_Y9_N0.coord_y = 9;
defparam asyncreset_ctrl_X17_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X17_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X18_Y10_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y10_SIG ));
defparam asyncreset_ctrl_X18_Y10_N0.coord_x = 25;
defparam asyncreset_ctrl_X18_Y10_N0.coord_y = 6;
defparam asyncreset_ctrl_X18_Y10_N0.coord_z = 0;
defparam asyncreset_ctrl_X18_Y10_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X18_Y11_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y11_SIG ));
defparam asyncreset_ctrl_X18_Y11_N0.coord_x = 25;
defparam asyncreset_ctrl_X18_Y11_N0.coord_y = 5;
defparam asyncreset_ctrl_X18_Y11_N0.coord_z = 0;
defparam asyncreset_ctrl_X18_Y11_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X18_Y13_N0(
	.Din(),
	.Dout(AsyncReset_X18_Y13_GND));
defparam asyncreset_ctrl_X18_Y13_N0.coord_x = 5;
defparam asyncreset_ctrl_X18_Y13_N0.coord_y = 17;
defparam asyncreset_ctrl_X18_Y13_N0.coord_z = 0;
defparam asyncreset_ctrl_X18_Y13_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X18_Y13_N1(
	.Din(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.Dout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q__AsyncReset_X18_Y13_INV ));
defparam asyncreset_ctrl_X18_Y13_N1.coord_x = 5;
defparam asyncreset_ctrl_X18_Y13_N1.coord_y = 17;
defparam asyncreset_ctrl_X18_Y13_N1.coord_z = 1;
defparam asyncreset_ctrl_X18_Y13_N1.AsyncCtrlMux = 2'b11;

alta_asyncctrl asyncreset_ctrl_X18_Y15_N0(
	.Din(),
	.Dout(AsyncReset_X18_Y15_GND));
defparam asyncreset_ctrl_X18_Y15_N0.coord_x = 6;
defparam asyncreset_ctrl_X18_Y15_N0.coord_y = 15;
defparam asyncreset_ctrl_X18_Y15_N0.coord_z = 0;
defparam asyncreset_ctrl_X18_Y15_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X18_Y16_N0(
	.Din(),
	.Dout(AsyncReset_X18_Y16_GND));
defparam asyncreset_ctrl_X18_Y16_N0.coord_x = 6;
defparam asyncreset_ctrl_X18_Y16_N0.coord_y = 17;
defparam asyncreset_ctrl_X18_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X18_Y16_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X18_Y16_N1(
	.Din(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.Dout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8]__AsyncReset_X18_Y16_SIG ));
defparam asyncreset_ctrl_X18_Y16_N1.coord_x = 6;
defparam asyncreset_ctrl_X18_Y16_N1.coord_y = 17;
defparam asyncreset_ctrl_X18_Y16_N1.coord_z = 1;
defparam asyncreset_ctrl_X18_Y16_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X18_Y17_N0(
	.Din(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.Dout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ));
defparam asyncreset_ctrl_X18_Y17_N0.coord_x = 5;
defparam asyncreset_ctrl_X18_Y17_N0.coord_y = 16;
defparam asyncreset_ctrl_X18_Y17_N0.coord_z = 0;
defparam asyncreset_ctrl_X18_Y17_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X18_Y18_N0(
	.Din(),
	.Dout(AsyncReset_X18_Y18_GND));
defparam asyncreset_ctrl_X18_Y18_N0.coord_x = 8;
defparam asyncreset_ctrl_X18_Y18_N0.coord_y = 16;
defparam asyncreset_ctrl_X18_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X18_Y18_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X18_Y19_N0(
	.Din(),
	.Dout(AsyncReset_X18_Y19_GND));
defparam asyncreset_ctrl_X18_Y19_N0.coord_x = 10;
defparam asyncreset_ctrl_X18_Y19_N0.coord_y = 15;
defparam asyncreset_ctrl_X18_Y19_N0.coord_z = 0;
defparam asyncreset_ctrl_X18_Y19_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X18_Y19_N1(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X18_Y19_SIG ));
defparam asyncreset_ctrl_X18_Y19_N1.coord_x = 10;
defparam asyncreset_ctrl_X18_Y19_N1.coord_y = 15;
defparam asyncreset_ctrl_X18_Y19_N1.coord_z = 1;
defparam asyncreset_ctrl_X18_Y19_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X18_Y20_N0(
	.Din(),
	.Dout(AsyncReset_X18_Y20_GND));
defparam asyncreset_ctrl_X18_Y20_N0.coord_x = 13;
defparam asyncreset_ctrl_X18_Y20_N0.coord_y = 16;
defparam asyncreset_ctrl_X18_Y20_N0.coord_z = 0;
defparam asyncreset_ctrl_X18_Y20_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X19_Y16_N0(
	.Din(),
	.Dout(AsyncReset_X19_Y16_GND));
defparam asyncreset_ctrl_X19_Y16_N0.coord_x = 4;
defparam asyncreset_ctrl_X19_Y16_N0.coord_y = 17;
defparam asyncreset_ctrl_X19_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X19_Y16_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X19_Y17_N0(
	.Din(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.Dout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ));
defparam asyncreset_ctrl_X19_Y17_N0.coord_x = 2;
defparam asyncreset_ctrl_X19_Y17_N0.coord_y = 15;
defparam asyncreset_ctrl_X19_Y17_N0.coord_z = 0;
defparam asyncreset_ctrl_X19_Y17_N0.AsyncCtrlMux = 2'b11;

alta_asyncctrl asyncreset_ctrl_X19_Y18_N0(
	.Din(),
	.Dout(AsyncReset_X19_Y18_GND));
defparam asyncreset_ctrl_X19_Y18_N0.coord_x = 7;
defparam asyncreset_ctrl_X19_Y18_N0.coord_y = 15;
defparam asyncreset_ctrl_X19_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X19_Y18_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X19_Y19_N0(
	.Din(),
	.Dout(AsyncReset_X19_Y19_GND));
defparam asyncreset_ctrl_X19_Y19_N0.coord_x = 9;
defparam asyncreset_ctrl_X19_Y19_N0.coord_y = 15;
defparam asyncreset_ctrl_X19_Y19_N0.coord_z = 0;
defparam asyncreset_ctrl_X19_Y19_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X19_Y8_N1(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X19_Y8_SIG ));
defparam asyncreset_ctrl_X19_Y8_N1.coord_x = 26;
defparam asyncreset_ctrl_X19_Y8_N1.coord_y = 6;
defparam asyncreset_ctrl_X19_Y8_N1.coord_z = 1;
defparam asyncreset_ctrl_X19_Y8_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X1_Y1_N0(
	.Din(\reset_init[5]~clkctrl_outclk ),
	.Dout(\reset_init[5]~clkctrl_outclk__AsyncReset_X1_Y1_INV ));
defparam asyncreset_ctrl_X1_Y1_N0.coord_x = 1;
defparam asyncreset_ctrl_X1_Y1_N0.coord_y = 12;
defparam asyncreset_ctrl_X1_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X1_Y1_N0.AsyncCtrlMux = 2'b11;

alta_asyncctrl asyncreset_ctrl_X1_Y7_N0(
	.Din(),
	.Dout(AsyncReset_X1_Y7_GND));
defparam asyncreset_ctrl_X1_Y7_N0.coord_x = 4;
defparam asyncreset_ctrl_X1_Y7_N0.coord_y = 11;
defparam asyncreset_ctrl_X1_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X1_Y7_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X21_Y14_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ));
defparam asyncreset_ctrl_X21_Y14_N0.coord_x = 21;
defparam asyncreset_ctrl_X21_Y14_N0.coord_y = 12;
defparam asyncreset_ctrl_X21_Y14_N0.coord_z = 0;
defparam asyncreset_ctrl_X21_Y14_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X21_Y15_N0(
	.Din(),
	.Dout(AsyncReset_X21_Y15_GND));
defparam asyncreset_ctrl_X21_Y15_N0.coord_x = 3;
defparam asyncreset_ctrl_X21_Y15_N0.coord_y = 15;
defparam asyncreset_ctrl_X21_Y15_N0.coord_z = 0;
defparam asyncreset_ctrl_X21_Y15_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X21_Y16_N0(
	.Din(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.Dout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X21_Y16_SIG ));
defparam asyncreset_ctrl_X21_Y16_N0.coord_x = 4;
defparam asyncreset_ctrl_X21_Y16_N0.coord_y = 15;
defparam asyncreset_ctrl_X21_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X21_Y16_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X21_Y17_N0(
	.Din(),
	.Dout(AsyncReset_X21_Y17_GND));
defparam asyncreset_ctrl_X21_Y17_N0.coord_x = 1;
defparam asyncreset_ctrl_X21_Y17_N0.coord_y = 15;
defparam asyncreset_ctrl_X21_Y17_N0.coord_z = 0;
defparam asyncreset_ctrl_X21_Y17_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X21_Y18_N0(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y18_SIG ));
defparam asyncreset_ctrl_X21_Y18_N0.coord_x = 9;
defparam asyncreset_ctrl_X21_Y18_N0.coord_y = 16;
defparam asyncreset_ctrl_X21_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X21_Y18_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X21_Y18_N1(
	.Din(),
	.Dout(AsyncReset_X21_Y18_GND));
defparam asyncreset_ctrl_X21_Y18_N1.coord_x = 9;
defparam asyncreset_ctrl_X21_Y18_N1.coord_y = 16;
defparam asyncreset_ctrl_X21_Y18_N1.coord_z = 1;
defparam asyncreset_ctrl_X21_Y18_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X21_Y19_N0(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ));
defparam asyncreset_ctrl_X21_Y19_N0.coord_x = 11;
defparam asyncreset_ctrl_X21_Y19_N0.coord_y = 15;
defparam asyncreset_ctrl_X21_Y19_N0.coord_z = 0;
defparam asyncreset_ctrl_X21_Y19_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X21_Y20_N0(
	.Din(),
	.Dout(AsyncReset_X21_Y20_GND));
defparam asyncreset_ctrl_X21_Y20_N0.coord_x = 10;
defparam asyncreset_ctrl_X21_Y20_N0.coord_y = 17;
defparam asyncreset_ctrl_X21_Y20_N0.coord_z = 0;
defparam asyncreset_ctrl_X21_Y20_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X22_Y14_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y14_SIG ));
defparam asyncreset_ctrl_X22_Y14_N0.coord_x = 21;
defparam asyncreset_ctrl_X22_Y14_N0.coord_y = 13;
defparam asyncreset_ctrl_X22_Y14_N0.coord_z = 0;
defparam asyncreset_ctrl_X22_Y14_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X22_Y14_N1(
	.Din(),
	.Dout(AsyncReset_X22_Y14_GND));
defparam asyncreset_ctrl_X22_Y14_N1.coord_x = 21;
defparam asyncreset_ctrl_X22_Y14_N1.coord_y = 13;
defparam asyncreset_ctrl_X22_Y14_N1.coord_z = 1;
defparam asyncreset_ctrl_X22_Y14_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X22_Y15_N0(
	.Din(),
	.Dout(AsyncReset_X22_Y15_GND));
defparam asyncreset_ctrl_X22_Y15_N0.coord_x = 21;
defparam asyncreset_ctrl_X22_Y15_N0.coord_y = 14;
defparam asyncreset_ctrl_X22_Y15_N0.coord_z = 0;
defparam asyncreset_ctrl_X22_Y15_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X22_Y15_N1(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y15_SIG ));
defparam asyncreset_ctrl_X22_Y15_N1.coord_x = 21;
defparam asyncreset_ctrl_X22_Y15_N1.coord_y = 14;
defparam asyncreset_ctrl_X22_Y15_N1.coord_z = 1;
defparam asyncreset_ctrl_X22_Y15_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X22_Y17_N0(
	.Din(),
	.Dout(AsyncReset_X22_Y17_GND));
defparam asyncreset_ctrl_X22_Y17_N0.coord_x = 5;
defparam asyncreset_ctrl_X22_Y17_N0.coord_y = 14;
defparam asyncreset_ctrl_X22_Y17_N0.coord_z = 0;
defparam asyncreset_ctrl_X22_Y17_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X22_Y18_N0(
	.Din(),
	.Dout(AsyncReset_X22_Y18_GND));
defparam asyncreset_ctrl_X22_Y18_N0.coord_x = 8;
defparam asyncreset_ctrl_X22_Y18_N0.coord_y = 15;
defparam asyncreset_ctrl_X22_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X22_Y18_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X22_Y19_N0(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X22_Y19_SIG ));
defparam asyncreset_ctrl_X22_Y19_N0.coord_x = 10;
defparam asyncreset_ctrl_X22_Y19_N0.coord_y = 16;
defparam asyncreset_ctrl_X22_Y19_N0.coord_z = 0;
defparam asyncreset_ctrl_X22_Y19_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X23_Y16_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ));
defparam asyncreset_ctrl_X23_Y16_N0.coord_x = 20;
defparam asyncreset_ctrl_X23_Y16_N0.coord_y = 10;
defparam asyncreset_ctrl_X23_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X23_Y16_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X23_Y19_N0(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X23_Y19_SIG ));
defparam asyncreset_ctrl_X23_Y19_N0.coord_x = 11;
defparam asyncreset_ctrl_X23_Y19_N0.coord_y = 16;
defparam asyncreset_ctrl_X23_Y19_N0.coord_z = 0;
defparam asyncreset_ctrl_X23_Y19_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X24_Y12_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y12_SIG ));
defparam asyncreset_ctrl_X24_Y12_N0.coord_x = 19;
defparam asyncreset_ctrl_X24_Y12_N0.coord_y = 10;
defparam asyncreset_ctrl_X24_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X24_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X24_Y15_N1(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ));
defparam asyncreset_ctrl_X24_Y15_N1.coord_x = 21;
defparam asyncreset_ctrl_X24_Y15_N1.coord_y = 10;
defparam asyncreset_ctrl_X24_Y15_N1.coord_z = 1;
defparam asyncreset_ctrl_X24_Y15_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X24_Y16_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ));
defparam asyncreset_ctrl_X24_Y16_N0.coord_x = 20;
defparam asyncreset_ctrl_X24_Y16_N0.coord_y = 12;
defparam asyncreset_ctrl_X24_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X24_Y16_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X24_Y18_N0(
	.Din(),
	.Dout(AsyncReset_X24_Y18_GND));
defparam asyncreset_ctrl_X24_Y18_N0.coord_x = 1;
defparam asyncreset_ctrl_X24_Y18_N0.coord_y = 11;
defparam asyncreset_ctrl_X24_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X24_Y18_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X24_Y19_N0(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ));
defparam asyncreset_ctrl_X24_Y19_N0.coord_x = 12;
defparam asyncreset_ctrl_X24_Y19_N0.coord_y = 16;
defparam asyncreset_ctrl_X24_Y19_N0.coord_z = 0;
defparam asyncreset_ctrl_X24_Y19_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X25_Y12_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y12_SIG ));
defparam asyncreset_ctrl_X25_Y12_N0.coord_x = 21;
defparam asyncreset_ctrl_X25_Y12_N0.coord_y = 9;
defparam asyncreset_ctrl_X25_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X25_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X25_Y13_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y13_SIG ));
defparam asyncreset_ctrl_X25_Y13_N0.coord_x = 22;
defparam asyncreset_ctrl_X25_Y13_N0.coord_y = 9;
defparam asyncreset_ctrl_X25_Y13_N0.coord_z = 0;
defparam asyncreset_ctrl_X25_Y13_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X25_Y15_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y15_SIG ));
defparam asyncreset_ctrl_X25_Y15_N0.coord_x = 20;
defparam asyncreset_ctrl_X25_Y15_N0.coord_y = 14;
defparam asyncreset_ctrl_X25_Y15_N0.coord_z = 0;
defparam asyncreset_ctrl_X25_Y15_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X25_Y15_N1(
	.Din(),
	.Dout(AsyncReset_X25_Y15_GND));
defparam asyncreset_ctrl_X25_Y15_N1.coord_x = 20;
defparam asyncreset_ctrl_X25_Y15_N1.coord_y = 14;
defparam asyncreset_ctrl_X25_Y15_N1.coord_z = 1;
defparam asyncreset_ctrl_X25_Y15_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X25_Y18_N0(
	.Din(),
	.Dout(AsyncReset_X25_Y18_GND));
defparam asyncreset_ctrl_X25_Y18_N0.coord_x = 2;
defparam asyncreset_ctrl_X25_Y18_N0.coord_y = 11;
defparam asyncreset_ctrl_X25_Y18_N0.coord_z = 0;
defparam asyncreset_ctrl_X25_Y18_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X25_Y19_N0(
	.Din(),
	.Dout(AsyncReset_X25_Y19_GND));
defparam asyncreset_ctrl_X25_Y19_N0.coord_x = 2;
defparam asyncreset_ctrl_X25_Y19_N0.coord_y = 12;
defparam asyncreset_ctrl_X25_Y19_N0.coord_z = 0;
defparam asyncreset_ctrl_X25_Y19_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X26_Y12_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y12_SIG ));
defparam asyncreset_ctrl_X26_Y12_N0.coord_x = 20;
defparam asyncreset_ctrl_X26_Y12_N0.coord_y = 9;
defparam asyncreset_ctrl_X26_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X26_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X26_Y13_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y13_SIG ));
defparam asyncreset_ctrl_X26_Y13_N0.coord_x = 22;
defparam asyncreset_ctrl_X26_Y13_N0.coord_y = 8;
defparam asyncreset_ctrl_X26_Y13_N0.coord_z = 0;
defparam asyncreset_ctrl_X26_Y13_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X26_Y15_N1(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ));
defparam asyncreset_ctrl_X26_Y15_N1.coord_x = 19;
defparam asyncreset_ctrl_X26_Y15_N1.coord_y = 14;
defparam asyncreset_ctrl_X26_Y15_N1.coord_z = 1;
defparam asyncreset_ctrl_X26_Y15_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X26_Y16_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y16_SIG ));
defparam asyncreset_ctrl_X26_Y16_N0.coord_x = 19;
defparam asyncreset_ctrl_X26_Y16_N0.coord_y = 12;
defparam asyncreset_ctrl_X26_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X26_Y16_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X28_Y9_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y9_SIG ));
defparam asyncreset_ctrl_X28_Y9_N0.coord_x = 24;
defparam asyncreset_ctrl_X28_Y9_N0.coord_y = 8;
defparam asyncreset_ctrl_X28_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X28_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X29_Y9_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ));
defparam asyncreset_ctrl_X29_Y9_N0.coord_x = 25;
defparam asyncreset_ctrl_X29_Y9_N0.coord_y = 8;
defparam asyncreset_ctrl_X29_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X29_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X2_Y7_N0(
	.Din(),
	.Dout(AsyncReset_X2_Y7_GND));
defparam asyncreset_ctrl_X2_Y7_N0.coord_x = 5;
defparam asyncreset_ctrl_X2_Y7_N0.coord_y = 11;
defparam asyncreset_ctrl_X2_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X2_Y7_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X33_Y12_N0(
	.Din(),
	.Dout(AsyncReset_X33_Y12_GND));
defparam asyncreset_ctrl_X33_Y12_N0.coord_x = 47;
defparam asyncreset_ctrl_X33_Y12_N0.coord_y = 15;
defparam asyncreset_ctrl_X33_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X33_Y12_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X33_Y16_N0(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ));
defparam asyncreset_ctrl_X33_Y16_N0.coord_x = 24;
defparam asyncreset_ctrl_X33_Y16_N0.coord_y = 9;
defparam asyncreset_ctrl_X33_Y16_N0.coord_z = 0;
defparam asyncreset_ctrl_X33_Y16_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X5_Y7_N1(
	.Din(),
	.Dout(AsyncReset_X5_Y7_GND));
defparam asyncreset_ctrl_X5_Y7_N1.coord_x = 8;
defparam asyncreset_ctrl_X5_Y7_N1.coord_y = 11;
defparam asyncreset_ctrl_X5_Y7_N1.coord_z = 1;
defparam asyncreset_ctrl_X5_Y7_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X9_Y7_N0(
	.Din(),
	.Dout(AsyncReset_X9_Y7_GND));
defparam asyncreset_ctrl_X9_Y7_N0.coord_x = 10;
defparam asyncreset_ctrl_X9_Y7_N0.coord_y = 11;
defparam asyncreset_ctrl_X9_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X9_Y7_N0.AsyncCtrlMux = 2'b00;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .coord_z = 13;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .mask = 16'h3000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X17_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .coord_z = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .coord_x = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .coord_z = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 (
	.A(vcc),
	.B(vcc),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .coord_z = 0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .mask = 16'h0FFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~24_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout_X18_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y16_GND),
	.SyncReset(SyncReset_X18_Y16_GND),
	.ShiftData(),
	.SyncLoad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout__SyncLoad_X18_Y16_SIG ),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .coord_z = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .mask = 16'hEE44;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~16 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.B(vcc),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~16_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~16 .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~16 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~16 .coord_z = 12;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~16 .mask = 16'hAA00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~16 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~16 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~16 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~16 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~16 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~16_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17 .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17 .coord_z = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17 .mask = 16'h8000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22_combout ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout_X18_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y16_GND),
	.SyncReset(SyncReset_X18_Y16_GND),
	.ShiftData(),
	.SyncLoad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout__SyncLoad_X18_Y16_SIG ),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .coord_z = 11;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .mask = 16'hDD88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout_X18_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y16_GND),
	.SyncReset(SyncReset_X18_Y16_GND),
	.ShiftData(),
	.SyncLoad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout__SyncLoad_X18_Y16_SIG ),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .coord_z = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .mask = 16'hDD88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~17_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.C(\altera_internal_jtag~TDIUTAP ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout_X18_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y16_GND),
	.SyncReset(SyncReset_X18_Y16_GND),
	.ShiftData(),
	.SyncLoad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout__SyncLoad_X18_Y16_SIG ),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .coord_z = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .mask = 16'hDD88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .coord_z = 0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .mask = 16'h2C27;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .coord_z = 13;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .mask = 16'h0A0D;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.B(vcc),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .coord_x = 8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .coord_z = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .mask = 16'hF0AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .coord_z = 14;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .mask = 16'h9384;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .coord_z = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .mask = 16'h0C8E;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .coord_z = 8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .mask = 16'h0436;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22 .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22 .coord_z = 9;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22 .mask = 16'h1E08;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~22 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23 .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23 .coord_z = 10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23 .mask = 16'h03D2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~24 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~23_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~24_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~24 .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~24 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~24 .coord_z = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~24 .mask = 16'h1F08;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~24 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~24 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~24 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~24 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~24 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.B(vcc),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .coord_z = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .mask = 16'hAAA0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .coord_z = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .mask = 16'hFFCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17_combout_X18_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .coord_z = 0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .mask = 16'hFF08;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17 .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17 .coord_z = 8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17 .mask = 16'hFEAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17_combout_X18_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .coord_z = 12;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .mask = 16'hAEEE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17_combout_X18_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~18_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .coord_z = 8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .mask = 16'h0CCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~15_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.D(\altera_internal_jtag~TDIUTAP ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17_combout_X17_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .coord_z = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .mask = 16'hDCCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .coord_z = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .mask = 16'h80F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .coord_z = 9;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .mask = 16'hCC0A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .coord_z = 14;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .mask = 16'hCC50;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .coord_z = 11;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .mask = 16'h44EF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~15 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~15_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~15 .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~15 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~15 .coord_z = 10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~15 .mask = 16'h0004;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~15 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~15 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~15 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~15 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~15 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .coord_z = 1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .mask = 16'h004C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .coord_z = 10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .mask = 16'h8000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .coord_z = 13;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .mask = 16'h0011;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .coord_z = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20_combout_X18_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y15_GND),
	.SyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13_combout__SyncReset_X18_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X18_Y15_GND),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~9_combout ),
	.Cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~10 ),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .coord_z = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .mask = 16'h55AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .CarryEnb = 1'b0;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13 .coord_z = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13 .mask = 16'hF2F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20 .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20 .coord_z = 13;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20 .mask = 16'hAEAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~10 ),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20_combout_X18_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y15_GND),
	.SyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13_combout__SyncReset_X18_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X18_Y15_GND),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~11_combout ),
	.Cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~12 ),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .coord_z = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .CarryEnb = 1'b0;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~12 ),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20_combout_X18_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y15_GND),
	.SyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13_combout__SyncReset_X18_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X18_Y15_GND),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~14_combout ),
	.Cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 ),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .coord_z = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .mask = 16'hA50A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .CarryEnb = 1'b0;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 ),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20_combout_X18_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y15_GND),
	.SyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13_combout__SyncReset_X18_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X18_Y15_GND),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~16_combout ),
	.Cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~17 ),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .coord_z = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .CarryEnb = 1'b0;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~17 ),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20_combout_X18_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y15_GND),
	.SyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13_combout__SyncReset_X18_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X18_Y15_GND),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~18_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .coord_z = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .mask = 16'hC3C3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.B(vcc),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout_X18_Y13_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y13_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .coord_z = 13;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .mask = 16'hFFAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.B(vcc),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout_X18_Y13_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y13_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .coord_z = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .mask = 16'h00AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.B(vcc),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout_X18_Y13_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y13_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .coord_z = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .mask = 16'hFFAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] (
	.A(\altera_internal_jtag~TDIUTAP ),
	.B(vcc),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout_X18_Y13_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y13_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .coord_z = 1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .mask = 16'h00AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y17_SIG_VCC ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X17_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .coord_z = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .mask = 16'h30B8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y17_SIG_VCC ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X17_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .coord_z = 12;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .mask = 16'hF078;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .coord_z = 9;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .mask = 16'h09A8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y13_SIG_VCC ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q__AsyncReset_X18_Y13_INV ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .coord_z = 8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .mask = 16'h7430;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .coord_z = 1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout_X19_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .coord_x = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .coord_z = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .mask = 16'hAAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .coord_z = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .mask = 16'h0080;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .coord_x = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .coord_z = 12;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .mask = 16'h3000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] (
	.A(),
	.B(),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.D(),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout_X19_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y16_GND),
	.SyncReset(SyncReset_X19_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y16_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .coord_x = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .coord_z = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .mask = 16'hFFFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout_X19_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .coord_x = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .coord_z = 11;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .mask = 16'hCCCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\altera_internal_jtag~TDIUTAP ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout_X19_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .coord_x = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .coord_z = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout_X19_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .coord_x = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .coord_z = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .mask = 16'hAAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .coord_x = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .coord_z = 0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .mask = 16'h0020;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout_X19_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .coord_x = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .coord_z = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .mask = 16'hAAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] (
	.A(),
	.B(),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.D(),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout_X19_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y16_GND),
	.SyncReset(SyncReset_X19_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y16_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .coord_x = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .coord_z = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .mask = 16'hFFFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout_X19_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .coord_x = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .coord_z = 14;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .mask = 16'hCCCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] (
	.A(),
	.B(),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.D(),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X17_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X17_Y17_SIG ),
	.SyncReset(SyncReset_X17_Y17_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X17_Y17_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .coord_z = 11;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .mask = 16'hFFFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .coord_z = 9;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .coord_z = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .mask = 16'hAAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] (
	.A(),
	.B(),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.D(),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(SyncReset_X18_Y17_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X18_Y17_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .coord_z = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .mask = 16'hFFFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] (
	.A(),
	.B(),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.D(),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X17_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X17_Y17_SIG ),
	.SyncReset(SyncReset_X17_Y17_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X17_Y17_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .coord_z = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .mask = 16'hFFFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X17_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X17_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .coord_z = 8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5] (
	.A(),
	.B(),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.D(),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5]~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(SyncReset_X18_Y17_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X18_Y17_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5]~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5] .coord_z = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5] .mask = 16'hFFFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [6]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6] .coord_z = 8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6] .mask = 16'hCCCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [7]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7] .coord_z = 9;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7] .mask = 16'hCCCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [8]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8]~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8]~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8] .coord_z = 14;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8] .mask = 16'hAAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [9]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9]~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9]~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9] .coord_z = 10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9] .mask = 16'hAAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~0_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .coord_z = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .mask = 16'hCCAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2 .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2 .coord_z = 14;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2 .mask = 16'hC0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[10] (
	.A(\altera_internal_jtag~TDIUTAP ),
	.B(vcc),
	.C(\~QIC_CREATED_GND~I_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q_X21_Y16_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X21_Y16_SIG ),
	.SyncReset(SyncReset_X21_Y16_GND),
	.ShiftData(),
	.SyncLoad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3]__SyncLoad_X21_Y16_SIG ),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~4_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[10] .coord_x = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[10] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[10] .coord_z = 11;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[10] .mask = 16'hAAF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[10] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[10] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[10] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[10] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[10] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .coord_z = 13;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .mask = 16'hCCF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~3_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .coord_z = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .mask = 16'hCCF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.B(vcc),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1 .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1 .coord_z = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1 .mask = 16'hF5A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~8_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~6_combout ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y17_SIG_VCC ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X17_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~9_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .coord_z = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .mask = 16'hF870;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~6 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~1_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~6_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~6 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~6 .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~6 .coord_z = 13;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~6 .mask = 16'hC0AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~6 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~6 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~6 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~6 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~6 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~7 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~7_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~7 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~7 .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~7 .coord_z = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~7 .mask = 16'hBB88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~7 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~7 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~7 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~7 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~7 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~8 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~7_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~8_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~8 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~8 .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~8 .coord_z = 1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~8 .mask = 16'hEEAE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~8 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~8 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~8 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~8 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~8 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~10_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .coord_z = 0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .mask = 16'hCCF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5]~q ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [6]),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~11_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .coord_z = 11;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .mask = 16'hAACC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[6] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [7]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~12_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [6]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[6] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[6] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[6] .coord_z = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[6] .mask = 16'hF0CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[6] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[6] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[6] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[6] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[6] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[7] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [8]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [7]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~13_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [7]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[7] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[7] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[7] .coord_z = 12;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[7] .mask = 16'hCCAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[7] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[7] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[7] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[7] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[7] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[8] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [9]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8]~q ),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [8]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~14_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [8]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[8] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[8] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[8] .coord_z = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[8] .mask = 16'hCCAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[8] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[8] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[8] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[8] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[8] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[9] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9]~q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [9]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout_X18_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X18_Y17_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~15_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [9]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[9] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[9] .coord_y = 16;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[9] .coord_z = 1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[9] .mask = 16'hCCF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[9] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[9] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[9] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[9] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[9] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11]_X19_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .coord_x = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .coord_z = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .mask = 16'h3333;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11]_X19_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .coord_x = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .coord_z = 14;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .mask = 16'hAAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11]_X19_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .coord_x = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .coord_z = 0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .mask = 16'h3333;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] (
	.A(),
	.B(),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.D(),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11]_X19_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ),
	.SyncReset(SyncReset_X19_Y17_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y17_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .coord_x = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .coord_z = 10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .mask = 16'hFFFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] (
	.A(),
	.B(),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.D(),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11]_X19_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ),
	.SyncReset(SyncReset_X19_Y17_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y17_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .coord_x = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .coord_z = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .mask = 16'hFFFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11]_X19_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ),
	.SyncReset(SyncReset_X19_Y17_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y17_VCC),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .coord_x = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .coord_z = 11;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .mask = 16'h0004;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11]_X19_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .coord_x = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .coord_z = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .mask = 16'hAAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] (
	.A(),
	.B(),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.D(),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11]_X19_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ),
	.SyncReset(SyncReset_X19_Y17_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y17_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .coord_x = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .coord_z = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .mask = 16'hFFFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] (
	.A(),
	.B(),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.D(),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11]_X19_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ),
	.SyncReset(SyncReset_X19_Y17_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y17_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .coord_x = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .coord_z = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .mask = 16'hFFFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.C(\altera_internal_jtag~TDIUTAP ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11]_X19_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ),
	.SyncReset(SyncReset_X19_Y17_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y17_VCC),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .coord_x = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .coord_z = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .mask = 16'h0001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout_X17_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y16_GND),
	.SyncReset(SyncReset_X17_Y16_GND),
	.ShiftData(),
	.SyncLoad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout__SyncLoad_X17_Y16_SIG ),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7_combout ),
	.Cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~8 ),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .coord_z = 1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .mask = 16'h55AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .CarryEnb = 1'b0;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~8 ),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout_X17_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y16_GND),
	.SyncReset(SyncReset_X17_Y16_GND),
	.ShiftData(),
	.SyncLoad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout__SyncLoad_X17_Y16_SIG ),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~11_combout ),
	.Cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~12 ),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .coord_z = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .mask = 16'hA505;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .CarryEnb = 1'b0;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~12 ),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout_X17_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y16_GND),
	.SyncReset(SyncReset_X17_Y16_GND),
	.ShiftData(),
	.SyncLoad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout__SyncLoad_X17_Y16_SIG ),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13_combout ),
	.Cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~14 ),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .coord_z = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .mask = 16'h5AAF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .CarryEnb = 1'b0;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~14 ),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout_X17_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y16_GND),
	.SyncReset(SyncReset_X17_Y16_GND),
	.ShiftData(),
	.SyncLoad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout__SyncLoad_X17_Y16_SIG ),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15_combout ),
	.Cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~16 ),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .coord_z = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .CarryEnb = 1'b0;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~16 ),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout_X17_Y16_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y16_GND),
	.SyncReset(SyncReset_X17_Y16_GND),
	.ShiftData(),
	.SyncLoad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout__SyncLoad_X17_Y16_SIG ),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .coord_z = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .mask = 16'h5A5A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .modeMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .coord_z = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .mask = 16'hEAC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 .coord_z = 9;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 .mask = 16'hCD05;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .coord_x = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .coord_z = 11;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .mask = 16'hFFFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y15_SIG_VCC ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q__AsyncReset_X17_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .coord_z = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .mask = 16'h88B8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 (
	.A(vcc),
	.B(vcc),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.D(\altera_internal_jtag~TMSUTAP ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .coord_z = 14;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 (
	.A(\altera_internal_jtag~TMSUTAP ),
	.B(\altera_internal_jtag~TDIUTAP ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .coord_z = 0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .mask = 16'hDF80;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.D(\altera_internal_jtag~TMSUTAP ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .coord_z = 1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .mask = 16'h0222;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .coord_z = 4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .mask = 16'hEE20;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.C(\altera_internal_jtag~TMSUTAP ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y13_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y13_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .coord_z = 14;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .mask = 16'hE000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.C(vcc),
	.D(\altera_internal_jtag~TMSUTAP ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X21_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .coord_x = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .coord_z = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .mask = 16'h10FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell (
	.A(vcc),
	.B(vcc),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .coord_x = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .coord_z = 12;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] (
	.A(vcc),
	.B(vcc),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.D(\altera_internal_jtag~TMSUTAP ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y17_SIG_VCC ),
	.AsyncReset(AsyncReset_X21_Y17_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .coord_x = 1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .coord_z = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .mask = 16'h00F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y17_SIG_VCC ),
	.AsyncReset(AsyncReset_X21_Y17_GND),
	.SyncReset(\altera_internal_jtag~TMSUTAP__SyncReset_X21_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X21_Y17_GND),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .coord_x = 1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .coord_z = 11;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .mask = 16'hFEFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.B(vcc),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.D(\altera_internal_jtag~TMSUTAP ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y17_SIG_VCC ),
	.AsyncReset(AsyncReset_X21_Y17_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .coord_x = 1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .coord_z = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .mask = 16'hFA00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y17_SIG_VCC ),
	.AsyncReset(AsyncReset_X21_Y17_GND),
	.SyncReset(\altera_internal_jtag~TMSUTAP__SyncReset_X21_Y17_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X21_Y17_GND),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .coord_x = 1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .coord_z = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .mask = 16'hFAFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.B(vcc),
	.C(vcc),
	.D(\altera_internal_jtag~TMSUTAP ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y17_SIG_VCC ),
	.AsyncReset(AsyncReset_X21_Y17_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .coord_x = 1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .coord_z = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .mask = 16'hAA00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.C(vcc),
	.D(\altera_internal_jtag~TMSUTAP ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y17_SIG_VCC ),
	.AsyncReset(AsyncReset_X21_Y17_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .coord_x = 1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .coord_z = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .mask = 16'hEE00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X17_Y15_GND),
	.SyncReset(\altera_internal_jtag~TMSUTAP__SyncReset_X17_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X17_Y15_GND),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .coord_z = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .mask = 16'hFFFB;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.C(\altera_internal_jtag~TMSUTAP ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X17_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .coord_z = 11;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .mask = 16'hF0E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] (
	.A(vcc),
	.B(vcc),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.D(\altera_internal_jtag~TMSUTAP ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X17_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .coord_z = 12;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .mask = 16'h00F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.B(vcc),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y13_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y13_GND),
	.SyncReset(\altera_internal_jtag~TMSUTAP__SyncReset_X18_Y13_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X18_Y13_GND),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .coord_z = 7;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .mask = 16'hFFFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.C(\altera_internal_jtag~TMSUTAP ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y13_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y13_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .coord_z = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y13_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y13_GND),
	.SyncReset(\altera_internal_jtag~TMSUTAP__SyncReset_X18_Y13_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X18_Y13_GND),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .coord_z = 12;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .mask = 16'hFAFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.C(\altera_internal_jtag~TMSUTAP ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y13_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y13_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .coord_z = 11;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.B(vcc),
	.C(\altera_internal_jtag~TMSUTAP ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y13_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y13_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .coord_z = 10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .mask = 16'hF0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] (
	.A(vcc),
	.B(vcc),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.D(\altera_internal_jtag~TMSUTAP ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X17_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .coord_z = 9;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\altera_internal_jtag~TMSUTAP ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X21_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .coord_x = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .coord_z = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X21_Y15_GND),
	.SyncReset(\altera_internal_jtag~TMSUTAP__SyncReset_X21_Y15_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X21_Y15_GND),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .coord_x = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .coord_z = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .mask = 16'h5A5A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X21_Y15_GND),
	.SyncReset(\altera_internal_jtag~TMSUTAP__SyncReset_X21_Y15_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X21_Y15_GND),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .coord_x = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .coord_z = 11;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .mask = 16'h7878;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .BypassEn = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout_X18_Y16_INV_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8]__AsyncReset_X18_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .coord_z = 14;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .mask = 16'h334F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.C(vcc),
	.D(\altera_internal_jtag~TDIUTAP ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y13_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y13_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .coord_x = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .coord_z = 0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .mask = 16'hFC30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .FeedbackMux = 1'b1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .coord_z = 8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .mask = 16'hF0CA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .coord_z = 10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .mask = 16'hD8D8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .coord_z = 12;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .mask = 16'hF0AC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .coord_z = 5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .mask = 16'hF0A2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .coord_x = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .coord_z = 6;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .mask = 16'hFCF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.Cout(),
	.Q());
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .coord_x = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .coord_y = 17;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .coord_z = 3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout_X19_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .coord_x = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .coord_z = 9;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .CarryEnb = 1'b1;

alta_slice \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.Cin(),
	.Qin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout_X19_Y17_SIG_SIG ),
	.AsyncReset(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]__AsyncReset_X19_Y17_INV ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.Cout(),
	.Q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ));
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .coord_x = 2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .coord_y = 15;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .coord_z = 8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .mask = 16'h1000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .modeMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .FeedbackMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .ShiftMux = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .BypassEn = 1'b0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .CarryEnb = 1'b1;

alta_slice \auto_hub|~GND (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_hub|~GND~combout ),
	.Cout(),
	.Q());
defparam \auto_hub|~GND .coord_x = 1;
defparam \auto_hub|~GND .coord_y = 1;
defparam \auto_hub|~GND .coord_z = 0;
defparam \auto_hub|~GND .mask = 16'h0000;
defparam \auto_hub|~GND .modeMux = 1'b0;
defparam \auto_hub|~GND .FeedbackMux = 1'b0;
defparam \auto_hub|~GND .ShiftMux = 1'b0;
defparam \auto_hub|~GND .BypassEn = 1'b0;
defparam \auto_hub|~GND .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_data_in_reg[0] (
	.A(vcc),
	.B(vcc),
	.C(\cam_data[0]~input_o ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_data_in_reg [0]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|acq_data_in_reg[0]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_data_in_reg [0]));
defparam \auto_signaltap_0|acq_data_in_reg[0] .coord_x = 17;
defparam \auto_signaltap_0|acq_data_in_reg[0] .coord_y = 15;
defparam \auto_signaltap_0|acq_data_in_reg[0] .coord_z = 8;
defparam \auto_signaltap_0|acq_data_in_reg[0] .mask = 16'hF0F0;
defparam \auto_signaltap_0|acq_data_in_reg[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_data_in_reg[1] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cam_data[1]~input_o ),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_data_in_reg [1]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|acq_data_in_reg[1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_data_in_reg [1]));
defparam \auto_signaltap_0|acq_data_in_reg[1] .coord_x = 17;
defparam \auto_signaltap_0|acq_data_in_reg[1] .coord_y = 15;
defparam \auto_signaltap_0|acq_data_in_reg[1] .coord_z = 11;
defparam \auto_signaltap_0|acq_data_in_reg[1] .mask = 16'hFF00;
defparam \auto_signaltap_0|acq_data_in_reg[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_data_in_reg[2] (
	.A(vcc),
	.B(vcc),
	.C(\cam_data[2]~input_o ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_data_in_reg [2]),
	.Clk(\clk~inputclkctrl_outclk_X13_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|acq_data_in_reg[2]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_data_in_reg [2]));
defparam \auto_signaltap_0|acq_data_in_reg[2] .coord_x = 17;
defparam \auto_signaltap_0|acq_data_in_reg[2] .coord_y = 14;
defparam \auto_signaltap_0|acq_data_in_reg[2] .coord_z = 8;
defparam \auto_signaltap_0|acq_data_in_reg[2] .mask = 16'hF0F0;
defparam \auto_signaltap_0|acq_data_in_reg[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_data_in_reg[3] (
	.A(),
	.B(),
	.C(\cam_data[3]~input_o ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_data_in_reg [3]),
	.Clk(\clk~inputclkctrl_outclk_X13_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y16_GND),
	.SyncReset(SyncReset_X13_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y16_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|acq_data_in_reg [3]));
defparam \auto_signaltap_0|acq_data_in_reg[3] .coord_x = 17;
defparam \auto_signaltap_0|acq_data_in_reg[3] .coord_y = 14;
defparam \auto_signaltap_0|acq_data_in_reg[3] .coord_z = 15;
defparam \auto_signaltap_0|acq_data_in_reg[3] .mask = 16'hFFFF;
defparam \auto_signaltap_0|acq_data_in_reg[3] .modeMux = 1'b1;
defparam \auto_signaltap_0|acq_data_in_reg[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[3] .BypassEn = 1'b1;
defparam \auto_signaltap_0|acq_data_in_reg[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_data_in_reg[4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cam_data[4]~input_o ),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_data_in_reg [4]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|acq_data_in_reg[4]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_data_in_reg [4]));
defparam \auto_signaltap_0|acq_data_in_reg[4] .coord_x = 17;
defparam \auto_signaltap_0|acq_data_in_reg[4] .coord_y = 15;
defparam \auto_signaltap_0|acq_data_in_reg[4] .coord_z = 3;
defparam \auto_signaltap_0|acq_data_in_reg[4] .mask = 16'hFF00;
defparam \auto_signaltap_0|acq_data_in_reg[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_data_in_reg[5] (
	.A(),
	.B(),
	.C(\cam_data[5]~input_o ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_data_in_reg [5]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(SyncReset_X12_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|acq_data_in_reg [5]));
defparam \auto_signaltap_0|acq_data_in_reg[5] .coord_x = 10;
defparam \auto_signaltap_0|acq_data_in_reg[5] .coord_y = 14;
defparam \auto_signaltap_0|acq_data_in_reg[5] .coord_z = 6;
defparam \auto_signaltap_0|acq_data_in_reg[5] .mask = 16'hFFFF;
defparam \auto_signaltap_0|acq_data_in_reg[5] .modeMux = 1'b1;
defparam \auto_signaltap_0|acq_data_in_reg[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[5] .BypassEn = 1'b1;
defparam \auto_signaltap_0|acq_data_in_reg[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_data_in_reg[6] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cam_data[6]~input_o ),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_data_in_reg [6]),
	.Clk(\clk~inputclkctrl_outclk_X11_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|acq_data_in_reg[6]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_data_in_reg [6]));
defparam \auto_signaltap_0|acq_data_in_reg[6] .coord_x = 16;
defparam \auto_signaltap_0|acq_data_in_reg[6] .coord_y = 15;
defparam \auto_signaltap_0|acq_data_in_reg[6] .coord_z = 11;
defparam \auto_signaltap_0|acq_data_in_reg[6] .mask = 16'hFF00;
defparam \auto_signaltap_0|acq_data_in_reg[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_data_in_reg[7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cam_data[7]~input_o ),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_data_in_reg [7]),
	.Clk(\clk~inputclkctrl_outclk_X11_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|acq_data_in_reg[7]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_data_in_reg [7]));
defparam \auto_signaltap_0|acq_data_in_reg[7] .coord_x = 16;
defparam \auto_signaltap_0|acq_data_in_reg[7] .coord_y = 15;
defparam \auto_signaltap_0|acq_data_in_reg[7] .coord_z = 8;
defparam \auto_signaltap_0|acq_data_in_reg[7] .mask = 16'hFF00;
defparam \auto_signaltap_0|acq_data_in_reg[7] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|acq_data_in_reg[7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_trigger_in_reg[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [0]),
	.C(\cam_data[0]~input_o ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [1]),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_trigger_in_reg [0]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(SyncReset_X12_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|p_match_out~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_trigger_in_reg [0]));
defparam \auto_signaltap_0|acq_trigger_in_reg[0] .coord_x = 10;
defparam \auto_signaltap_0|acq_trigger_in_reg[0] .coord_y = 14;
defparam \auto_signaltap_0|acq_trigger_in_reg[0] .coord_z = 7;
defparam \auto_signaltap_0|acq_trigger_in_reg[0] .mask = 16'hFC1D;
defparam \auto_signaltap_0|acq_trigger_in_reg[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[0] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[0] .BypassEn = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_trigger_in_reg[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [3]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [5]),
	.C(\cam_data[1]~input_o ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [4]),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_trigger_in_reg [1]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y18_GND),
	.SyncReset(SyncReset_X12_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y18_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|p_match_out~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_trigger_in_reg [1]));
defparam \auto_signaltap_0|acq_trigger_in_reg[1] .coord_x = 11;
defparam \auto_signaltap_0|acq_trigger_in_reg[1] .coord_y = 14;
defparam \auto_signaltap_0|acq_trigger_in_reg[1] .coord_z = 3;
defparam \auto_signaltap_0|acq_trigger_in_reg[1] .mask = 16'hFA1B;
defparam \auto_signaltap_0|acq_trigger_in_reg[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[1] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[1] .BypassEn = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_trigger_in_reg[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [6]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [7]),
	.C(\cam_data[2]~input_o ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [8]),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_trigger_in_reg [2]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y18_GND),
	.SyncReset(SyncReset_X12_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y18_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|p_match_out~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_trigger_in_reg [2]));
defparam \auto_signaltap_0|acq_trigger_in_reg[2] .coord_x = 11;
defparam \auto_signaltap_0|acq_trigger_in_reg[2] .coord_y = 14;
defparam \auto_signaltap_0|acq_trigger_in_reg[2] .coord_z = 12;
defparam \auto_signaltap_0|acq_trigger_in_reg[2] .mask = 16'hCADB;
defparam \auto_signaltap_0|acq_trigger_in_reg[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[2] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[2] .BypassEn = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_trigger_in_reg[3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [9]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [10]),
	.C(\cam_data[3]~input_o ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [11]),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_trigger_in_reg [3]),
	.Clk(\clk~inputclkctrl_outclk_X13_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y18_GND),
	.SyncReset(SyncReset_X13_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y18_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|p_match_out~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_trigger_in_reg [3]));
defparam \auto_signaltap_0|acq_trigger_in_reg[3] .coord_x = 10;
defparam \auto_signaltap_0|acq_trigger_in_reg[3] .coord_y = 12;
defparam \auto_signaltap_0|acq_trigger_in_reg[3] .coord_z = 11;
defparam \auto_signaltap_0|acq_trigger_in_reg[3] .mask = 16'hCADB;
defparam \auto_signaltap_0|acq_trigger_in_reg[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[3] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[3] .BypassEn = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_trigger_in_reg[4] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [12]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [13]),
	.C(\cam_data[4]~input_o ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [14]),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_trigger_in_reg [4]),
	.Clk(\clk~inputclkctrl_outclk_X13_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y18_GND),
	.SyncReset(SyncReset_X13_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y18_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|p_match_out~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_trigger_in_reg [4]));
defparam \auto_signaltap_0|acq_trigger_in_reg[4] .coord_x = 10;
defparam \auto_signaltap_0|acq_trigger_in_reg[4] .coord_y = 12;
defparam \auto_signaltap_0|acq_trigger_in_reg[4] .coord_z = 9;
defparam \auto_signaltap_0|acq_trigger_in_reg[4] .mask = 16'hCADB;
defparam \auto_signaltap_0|acq_trigger_in_reg[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[4] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[4] .BypassEn = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_trigger_in_reg[5] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [16]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [15]),
	.C(\cam_data[5]~input_o ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [17]),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_trigger_in_reg [5]),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(SyncReset_X12_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|p_match_out~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_trigger_in_reg [5]));
defparam \auto_signaltap_0|acq_trigger_in_reg[5] .coord_x = 10;
defparam \auto_signaltap_0|acq_trigger_in_reg[5] .coord_y = 14;
defparam \auto_signaltap_0|acq_trigger_in_reg[5] .coord_z = 3;
defparam \auto_signaltap_0|acq_trigger_in_reg[5] .mask = 16'hACBD;
defparam \auto_signaltap_0|acq_trigger_in_reg[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[5] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[5] .BypassEn = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_trigger_in_reg[6] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [19]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [20]),
	.C(\cam_data[6]~input_o ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [18]),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_trigger_in_reg [6]),
	.Clk(\clk~inputclkctrl_outclk_X11_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y14_GND),
	.SyncReset(SyncReset_X11_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y14_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|p_match_out~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_trigger_in_reg [6]));
defparam \auto_signaltap_0|acq_trigger_in_reg[6] .coord_x = 9;
defparam \auto_signaltap_0|acq_trigger_in_reg[6] .coord_y = 14;
defparam \auto_signaltap_0|acq_trigger_in_reg[6] .coord_z = 2;
defparam \auto_signaltap_0|acq_trigger_in_reg[6] .mask = 16'hAFB1;
defparam \auto_signaltap_0|acq_trigger_in_reg[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[6] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[6] .BypassEn = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|acq_trigger_in_reg[7] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [21]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [22]),
	.C(\cam_data[7]~input_o ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [23]),
	.Cin(),
	.Qin(\auto_signaltap_0|acq_trigger_in_reg [7]),
	.Clk(\clk~inputclkctrl_outclk_X11_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y14_GND),
	.SyncReset(SyncReset_X11_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y14_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|p_match_out~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|acq_trigger_in_reg [7]));
defparam \auto_signaltap_0|acq_trigger_in_reg[7] .coord_x = 9;
defparam \auto_signaltap_0|acq_trigger_in_reg[7] .coord_y = 14;
defparam \auto_signaltap_0|acq_trigger_in_reg[7] .coord_z = 7;
defparam \auto_signaltap_0|acq_trigger_in_reg[7] .mask = 16'hCADB;
defparam \auto_signaltap_0|acq_trigger_in_reg[7] .modeMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[7] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|acq_trigger_in_reg[7] .BypassEn = 1'b1;
defparam \auto_signaltap_0|acq_trigger_in_reg[7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [3]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [0]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~0 .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~0 .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~0 .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~0 .mask = 16'h0001;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~1 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [6]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [5]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [4]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~1_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~1 .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~1 .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~1 .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~1 .mask = 16'h0001;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~1 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~1 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~1 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~1 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~1 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~2 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [10]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [11]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [9]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [8]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~2_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~2 .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~2 .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~2 .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~2 .mask = 16'h0001;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~2 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~2 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~2 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~2 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~2 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~3 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [15]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [13]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [12]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [14]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~3_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~3 .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~3 .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~3 .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~3 .mask = 16'h0001;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~3 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~3 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~3 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~3 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~3 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~0_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~1_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~3_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4 .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4 .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4 .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4 .mask = 16'h8000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~5 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [19]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [18]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [16]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [17]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~5_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~5 .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~5 .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~5 .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~5 .mask = 16'h0001;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~5 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~5 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~5 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~5 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~5 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~6 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [23]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [22]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [21]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [20]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~6_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~6 .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~6 .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~6 .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~6 .mask = 16'h0001;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~6 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~6 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~6 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~6 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~6 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~7 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [27]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [26]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [25]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [24]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~7_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~7 .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~7 .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~7 .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~7 .mask = 16'h0001;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~7 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~7 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~7 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~7 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~7 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~8 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [30]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [31]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [28]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [29]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~8_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~8 .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~8 .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~8 .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~8 .mask = 16'h0001;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~8 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~8 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~8 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~8 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~8 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~7_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~6_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~8_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9 .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9 .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9 .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9 .mask = 16'h8000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0] (
	.A(vcc),
	.B(\auto_signaltap_0|acq_data_in_reg [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1] (
	.A(\auto_signaltap_0|acq_data_in_reg [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2] (
	.A(vcc),
	.B(\auto_signaltap_0|acq_data_in_reg [2]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2]~q ),
	.Clk(\clk~inputclkctrl_outclk_X13_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3] (
	.A(\auto_signaltap_0|acq_data_in_reg [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3]~q ),
	.Clk(\clk~inputclkctrl_outclk_X13_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|acq_data_in_reg [4]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(SyncReset_X12_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y16_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5] (
	.A(\auto_signaltap_0|acq_data_in_reg [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6] (
	.A(\auto_signaltap_0|acq_data_in_reg [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6]~q ),
	.Clk(\clk~inputclkctrl_outclk_X11_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6] .coord_x = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7] (
	.A(vcc),
	.B(\auto_signaltap_0|acq_data_in_reg [7]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7]~q ),
	.Clk(\clk~inputclkctrl_outclk_X11_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7] .coord_x = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][1]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][2]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2]~q ),
	.Clk(\clk~inputclkctrl_outclk_X13_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][3]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3]~q ),
	.Clk(\clk~inputclkctrl_outclk_X13_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][4]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][5]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][6]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6]~q ),
	.Clk(\clk~inputclkctrl_outclk_X11_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6] .coord_x = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[0][7]~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7]~q ),
	.Clk(\clk~inputclkctrl_outclk_X11_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y16_GND),
	.SyncReset(SyncReset_X11_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y16_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7] .coord_x = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][0]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][1]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][2]~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2]~q ),
	.Clk(\clk~inputclkctrl_outclk_X13_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y16_GND),
	.SyncReset(SyncReset_X13_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y16_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][3]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3]~q ),
	.Clk(\clk~inputclkctrl_outclk_X13_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][4]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][5]~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(SyncReset_X12_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][6]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6]~q ),
	.Clk(\clk~inputclkctrl_outclk_X11_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6] .coord_x = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[1][7]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7]~q ),
	.Clk(\clk~inputclkctrl_outclk_X11_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7] .coord_x = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][0]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][1]~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(SyncReset_X12_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y16_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][2]~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2]~q ),
	.Clk(\clk~inputclkctrl_outclk_X13_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y16_GND),
	.SyncReset(SyncReset_X13_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y16_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][3]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3]~q ),
	.Clk(\clk~inputclkctrl_outclk_X13_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][4]~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y16_GND),
	.SyncReset(SyncReset_X12_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y16_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][5]~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5]~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(SyncReset_X12_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][6]~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6]~q ),
	.Clk(\clk~inputclkctrl_outclk_X11_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y16_GND),
	.SyncReset(SyncReset_X11_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y16_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6] .coord_x = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[2][7]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7]~q ),
	.Clk(\clk~inputclkctrl_outclk_X11_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7] .coord_x = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [0]),
	.Clk(\clk~inputclkctrl_outclk_X14_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X14_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[0]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[0] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[0] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[0] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[0] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[1] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [1]),
	.Clk(\clk~inputclkctrl_outclk_X14_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X14_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[1] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[1] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[1] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[2] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [2]),
	.Clk(\clk~inputclkctrl_outclk_X14_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X14_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[2]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[2] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[2] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[2] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[2] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[3] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3]~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [3]),
	.Clk(\clk~inputclkctrl_outclk_X14_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X14_Y16_GND),
	.SyncReset(SyncReset_X14_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y16_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[3] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[3] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[3] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[3] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[3] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[3] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[4] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [4]),
	.Clk(\clk~inputclkctrl_outclk_X14_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X14_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[4]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[4] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[4] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[4] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[5] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [5]),
	.Clk(\clk~inputclkctrl_outclk_X14_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X14_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[5]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[5] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[5] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[5] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[5] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[6] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [6]),
	.Clk(\clk~inputclkctrl_outclk_X14_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X14_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[6]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[6] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[6] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[6] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[6] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed~q ),
	.Clk(\clk~inputclkctrl_outclk_X21_Y20_SIG_VCC ),
	.AsyncReset(AsyncReset_X21_Y20_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed .coord_y = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed .mask = 16'h00FF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out (
	.A(\altera_internal_jtag~TDIUTAP ),
	.B(vcc),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y18_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out .mask = 16'hAAF0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0 (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0 .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0 .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0 .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0 .mask = 16'h0C00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [0]),
	.Clk(\clk~inputclkctrl_outclk_X18_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[0]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[0] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[0] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[0] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[1] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [1]),
	.Clk(\clk~inputclkctrl_outclk_X18_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[1] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[1] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[1] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [2]),
	.Clk(\clk~inputclkctrl_outclk_X18_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[2]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[2] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[2] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[2] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[2] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run~q ),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [2]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [3]),
	.Clk(\clk~inputclkctrl_outclk_X18_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y19_GND),
	.SyncReset(SyncReset_X18_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X18_Y19_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[3] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[3] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[3] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[3] .mask = 16'hA0A0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[3] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[3] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|Add0~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [3]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [1]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|Add0~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|Add0~0 .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|Add0~0 .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|Add0~0 .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|Add0~0 .mask = 16'h6CCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|Add0~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|Add0~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|Add0~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|Add0~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|Add0~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [1]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~3_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12_combout_X22_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y17_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~4_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[0] .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[0] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[0] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[0] .mask = 16'h00F8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~6_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [2]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal~combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12_combout_X22_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y17_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~7_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[1] .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[1] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[1] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[1] .mask = 16'h0E0A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [3]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal~combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~8_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12_combout_X22_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y17_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~9_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2] .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2] .mask = 16'h0F08;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12 (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12 .coord_x = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12 .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12 .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12 .mask = 16'hFCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal~combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~10_combout ),
	.C(\altera_internal_jtag~TDIUTAP ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12_combout_X22_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y17_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~11_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[3] .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[3] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[3] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[3] .mask = 16'h5444;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~10 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [0]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [1]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~10_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~10 .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~10 .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~10 .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~10 .mask = 16'h5E00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~10 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~10 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~10 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~10 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~10 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2 (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [3]),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2 .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2 .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2 .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2 .mask = 16'h0033;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~3 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [0]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [1]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~3_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~3 .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~3 .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~3 .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~3 .mask = 16'h6E00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~3 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~3 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~3 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~3 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~3 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~5 (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [1]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~5_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~5 .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~5 .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~5 .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~5 .mask = 16'h0FFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~5 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~5 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~5 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~5 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~5 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~6 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [3]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [1]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~6_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~6 .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~6 .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~6 .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~6 .mask = 16'h0031;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~6 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~6 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~6 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~6 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~6 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~8 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [0]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [1]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~8_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~8 .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~8 .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~8 .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~8 .mask = 16'h6500;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~8 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~8 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~8 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~8 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~8 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal (
	.A(vcc),
	.B(vcc),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal~combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal .coord_x = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal .mask = 16'hF000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10_combout_X22_Y17_SIG_INV ),
	.AsyncReset(AsyncReset_X22_Y17_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter~11_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[0] .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[0] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[0] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[0] .mask = 16'h020A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[0] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal~combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [0]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10_combout_X22_Y17_SIG_INV ),
	.AsyncReset(AsyncReset_X22_Y17_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter~8_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[1] .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[1] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[1] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[1] .mask = 16'h1400;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[1] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR~5_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|clear_signal~combout ),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10_combout_X22_Y17_SIG_INV ),
	.AsyncReset(AsyncReset_X22_Y17_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter~7_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[2] .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[2] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[2] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[2] .mask = 16'h2100;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[2] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|Add0~0_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10_combout_X22_Y17_SIG_INV ),
	.AsyncReset(AsyncReset_X22_Y17_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter~9_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3] .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3] .mask = 16'h20A0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10 .coord_x = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10 .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10 .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10 .mask = 16'h45CF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [3]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [1]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6 .coord_x = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6 .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6 .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6 .mask = 16'hFFFB;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~6 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0]~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed [0]),
	.Clk(\clk~inputclkctrl_outclk_X21_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X21_Y18_GND),
	.SyncReset(SyncReset_X21_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X21_Y18_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed[0] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed[0] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed[0] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed[0] .mask = 16'h0A08;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed[0] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed[0] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[0] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [1]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[0]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[0] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[0] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[0] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[0] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[10] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [11]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [10]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X13_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X13_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[10]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [10]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[10] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[10] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[10] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[10] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[10] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[10] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[10] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[10] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[10] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[11] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [12]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [11]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X13_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X13_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[11]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [11]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[11] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[11] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[11] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[11] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[11] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[11] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[11] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[11] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[11] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[12] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [13]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [12]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X13_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X13_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[12]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [12]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[12] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[12] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[12] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[12] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[12] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[12] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[12] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[12] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[12] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[13] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [14]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [13]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X13_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X13_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[13]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [13]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[13] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[13] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[13] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[13] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[13] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[13] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[13] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[13] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[13] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[14] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [15]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [14]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X13_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X13_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[14]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [14]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[14] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[14] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[14] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[14] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[14] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[14] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[14] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[14] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[14] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[15] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [16]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [15]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X11_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X11_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[15]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [15]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[15] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[15] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[15] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[15] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[15] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[15] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[15] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[15] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[15] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[16] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [17]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [16]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X11_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X11_Y14_SIG ),
	.SyncReset(SyncReset_X11_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y14_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [16]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[16] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[16] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[16] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[16] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[16] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[16] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[16] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[16] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[16] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[17] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [18]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [17]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X11_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X11_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[17]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [17]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[17] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[17] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[17] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[17] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[17] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[17] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[17] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[17] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[17] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[18] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [19]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [18]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X11_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X11_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[18]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [18]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[18] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[18] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[18] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[18] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[18] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[18] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[18] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[18] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[18] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[19] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [20]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [19]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X11_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X11_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[19]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [19]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[19] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[19] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[19] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[19] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[19] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[19] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[19] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[19] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[19] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [2]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[1] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[1] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[1] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[1] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[20] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [21]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [20]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X11_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X11_Y14_SIG ),
	.SyncReset(SyncReset_X11_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y14_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [20]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[20] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[20] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[20] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[20] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[20] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[20] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[20] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[20] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[20] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[21] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [22]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [21]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X11_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X11_Y14_SIG ),
	.SyncReset(SyncReset_X11_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y14_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [21]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[21] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[21] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[21] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[21] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[21] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[21] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[21] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[21] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[21] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[22] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [23]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [22]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X11_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X11_Y14_SIG ),
	.SyncReset(SyncReset_X11_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y14_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [22]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[22] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[22] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[22] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[22] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[22] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[22] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[22] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[22] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[22] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[23] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\altera_internal_jtag~TDIUTAP ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [23]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X11_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X11_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[23]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [23]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[23] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[23] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[23] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[23] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[23] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[23] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[23] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[23] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[23] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[2]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[2] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[2] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[2] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[2] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[3] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [4]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y18_SIG ),
	.SyncReset(SyncReset_X12_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y18_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[3] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[3] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[3] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[3] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[3] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[3] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[4] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [5]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y18_SIG ),
	.SyncReset(SyncReset_X12_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y18_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[4] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[4] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[4] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[4] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[4] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[4] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[5] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[5]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[5] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[5] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[5] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[5] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[6] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [7]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[6]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[6] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[6] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[6] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[6] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [8]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [7]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[7]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [7]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[7] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[7] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[7] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[7] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[8] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [9]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [8]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[8]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [8]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[8] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[8] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[8] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[8] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[8] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[8] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[8] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[8] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[8] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[9] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [10]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [9]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X13_Y18_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X13_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[9]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [9]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[9] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[9] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[9] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[9] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[9] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[9] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[9] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[9] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs[9] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff (
	.A(vcc),
	.B(\auto_signaltap_0|acq_trigger_in_reg [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|holdff~q ),
	.B(\auto_signaltap_0|acq_trigger_in_reg [0]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|p_match_out~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [2]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|p_match_out~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff .mask = 16'h60F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff (
	.A(),
	.B(),
	.C(\auto_signaltap_0|acq_trigger_in_reg [1]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y18_GND),
	.SyncReset(SyncReset_X12_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y18_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|holdff~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [5]),
	.C(\auto_signaltap_0|acq_trigger_in_reg [1]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|p_match_out~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|p_match_out~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff .mask = 16'h7B00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff (
	.A(vcc),
	.B(\auto_signaltap_0|acq_trigger_in_reg [2]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|holdff~q ),
	.B(\auto_signaltap_0|acq_trigger_in_reg [2]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|p_match_out~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [8]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|p_match_out~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff .mask = 16'h60F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff (
	.A(\auto_signaltap_0|acq_trigger_in_reg [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff~q ),
	.Clk(\clk~inputclkctrl_outclk_X13_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff (
	.A(\auto_signaltap_0|acq_trigger_in_reg [3]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|holdff~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|p_match_out~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [11]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff~q ),
	.Clk(\clk~inputclkctrl_outclk_X13_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|p_match_out~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff .mask = 16'h60F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff (
	.A(),
	.B(),
	.C(\auto_signaltap_0|acq_trigger_in_reg [4]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff~q ),
	.Clk(\clk~inputclkctrl_outclk_X13_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y18_GND),
	.SyncReset(SyncReset_X13_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y18_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [14]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|holdff~q ),
	.C(\auto_signaltap_0|acq_trigger_in_reg [4]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|p_match_out~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff~q ),
	.Clk(\clk~inputclkctrl_outclk_X13_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X13_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|p_match_out~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff .mask = 16'h7D00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff (
	.A(\auto_signaltap_0|acq_trigger_in_reg [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff (
	.A(\auto_signaltap_0|acq_trigger_in_reg [5]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|holdff~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [17]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|p_match_out~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff~q ),
	.Clk(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X12_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|p_match_out~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff .mask = 16'h6F00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff (
	.A(vcc),
	.B(\auto_signaltap_0|acq_trigger_in_reg [6]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff~q ),
	.Clk(\clk~inputclkctrl_outclk_X11_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|holdff~q ),
	.B(\auto_signaltap_0|acq_trigger_in_reg [6]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|p_match_out~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [20]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff~q ),
	.Clk(\clk~inputclkctrl_outclk_X11_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|p_match_out~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff .mask = 16'h60F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff (
	.A(),
	.B(),
	.C(\auto_signaltap_0|acq_trigger_in_reg [7]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff~q ),
	.Clk(\clk~inputclkctrl_outclk_X11_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y14_GND),
	.SyncReset(SyncReset_X11_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y14_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff (
	.A(\auto_signaltap_0|acq_trigger_in_reg [7]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|holdff~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|p_match_out~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [23]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff~q ),
	.Clk(\clk~inputclkctrl_outclk_X11_Y14_SIG_VCC ),
	.AsyncReset(AsyncReset_X11_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|p_match_out~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff .mask = 16'h60F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~1_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run~q ),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~q ),
	.Clk(\clk~inputclkctrl_outclk_X18_Y19_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X18_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~2_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed .mask = 16'hB830;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:4:sm1|regoutff~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:3:sm1|regoutff~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:2:sm1|regoutff~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:1:sm1|regoutff~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~0 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~0 .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~0 .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~0 .mask = 16'h8000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~1 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:0:sm1|regoutff~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:5:sm1|regoutff~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:7:sm1|regoutff~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_modules_gen:0:trigger_match|gen_sbpmg_pipeline_less_than_two:sm0:6:sm1|regoutff~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~1_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~1 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~1 .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~1 .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~1 .mask = 16'h8000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~1 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~1 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~1 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~1 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~1 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [1]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(SyncReset_X21_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X21_Y19_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter~6_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[0] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[0] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[0] .mask = 16'h0032;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[0] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[0] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [2]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[1] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[1] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[1] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[2] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [3]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(SyncReset_X21_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X21_Y19_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[2] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[2] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[2] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[2] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[2] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[2] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [4]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[3]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[3] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[3] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[3] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[3] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[4] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [5]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(SyncReset_X21_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X21_Y19_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[4] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[4] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[4] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[4] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[4] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[5] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [6]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(SyncReset_X21_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X21_Y19_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[5] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[5] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[5] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[5] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[5] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[5] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[6] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [7]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[6]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[6] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[6] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[6] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[7] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [8]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [7]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[7]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [7]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[7] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[7] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[7] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[7] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[8] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [9]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [8]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[8]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [8]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[8] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[8] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[8] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[8] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[8] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[8] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[8] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[8] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[8] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[9] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|basic_multi_level_mbpm_trigger_gen:multi_level_mbpm|trigger_condition_deserialize|dffs [0]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [9]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X12_Y14_SIG ),
	.SyncReset(SyncReset_X12_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X12_Y14_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [9]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[9] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[9] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[9] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[9] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[9] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[9] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[9] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[9] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs[9] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [3]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run~q ),
	.Clk(\clk~inputclkctrl_outclk_X18_Y19_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X18_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run .mask = 16'hD555;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|run .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[0]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[0] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[0] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[0] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[1] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [2]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[1] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[1] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[1] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[2] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [3]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(SyncReset_X21_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X21_Y19_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[2] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[2] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[2] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[2] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[2] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[2] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[3] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[3]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[3] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[3] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[3] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[3] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[0] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0]~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [0]),
	.Clk(\clk~inputclkctrl_outclk_X14_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X14_Y18_GND),
	.SyncReset(SyncReset_X14_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y18_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[0] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[0] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[0] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[0] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[0] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[0] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[1] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [1]),
	.Clk(\clk~inputclkctrl_outclk_X14_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X14_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[1] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[1] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[1] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[1] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[2] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2]~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [2]),
	.Clk(\clk~inputclkctrl_outclk_X14_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X14_Y18_GND),
	.SyncReset(SyncReset_X14_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y18_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[2] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[2] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[2] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[2] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[2] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[2] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[3] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [3]),
	.Clk(\clk~inputclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[3]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[3] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[3] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[3] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[3] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[4] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4]~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [4]),
	.Clk(\clk~inputclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y16_GND),
	.SyncReset(SyncReset_X16_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y16_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[4] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[4] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[4] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[4] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[4] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [5]),
	.Clk(\clk~inputclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[5]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[5] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[5] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[5] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[5] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[6] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [6]),
	.Clk(\clk~inputclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y16_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[6]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[6] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[6] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[6] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~q ),
	.Clk(\clk~inputclkctrl_outclk_X18_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg .mask = 16'hFFF0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run~q ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~0 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~0 .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~0 .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~0 .mask = 16'hAAA8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8]~q ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0 .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0 .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0 .mask = 16'h2000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8]~q ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1 .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1 .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1 .mask = 16'h2000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2 (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [0]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2 .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2 .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2 .mask = 16'hFFCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~q ),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all .mask = 16'hFFC0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all .CarryEnb = 1'b1;

alta_io_gclk \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl (
	.inclk(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~q ),
	.outclk(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl .coord_x = 49;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl .coord_z = 2;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~q ),
	.B(vcc),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run~q ),
	.Clk(\clk~inputclkctrl_outclk_X18_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run .mask = 16'hFF55;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr .mask = 16'hFF3F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [0]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [1]),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X24_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ),
	.SyncReset(SyncReset_X24_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X24_Y19_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[0] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[0] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[0] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[0] .mask = 16'hE2C0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[0] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[0] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [2]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X24_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[1] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[1] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[1] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[1] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X24_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[2]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[2] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[2] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[2] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[2] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[3] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [4]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X24_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[3]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[3] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[3] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[3] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[3] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[4] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [5]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X24_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[4]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[4] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[4] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[4] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[4] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[5] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[5]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[5] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[5] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[5] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[5] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[6] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[6]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[6] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[6] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[6] .mask = 16'hAAAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped~q ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed~q ),
	.Clk(\clk~inputclkctrl_outclk_X18_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~0_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~1 ),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~0 .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~0 .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~0 .mask = 16'h55AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~0 .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~11 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [4]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~11_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~12 ),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~11 .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~11 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~11 .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~11 .mask = 16'hA50A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~11 .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~11 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~11 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~11 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~11 .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~14 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~12 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~14_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~15 ),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~14 .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~14 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~14 .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~14 .mask = 16'h5A5F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~14 .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~14 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~14 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~14 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~14 .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~17 (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [6]),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~17_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~18 ),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~17 .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~17 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~17 .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~17 .mask = 16'hC30C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~17 .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~17 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~17 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~17 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~17 .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~2 (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~2_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~3 ),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~2 .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~2 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~2 .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~2 .mask = 16'h3C3F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~2 .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~2 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~2 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~2 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~2 .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~20 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [7]),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~18 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~20_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~20 .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~20 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~20 .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~20 .mask = 16'h0FF0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~20 .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~20 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~20 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~20 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~20 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~5 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [2]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~5_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~6 ),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~5 .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~5 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~5 .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~5 .mask = 16'hA50A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~5 .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~5 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~5 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~5 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~5 .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~8 (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~6 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~8_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~9 ),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~8 .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~8 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~8 .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~8 .mask = 16'h3C3F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~8 .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~8 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~8 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~8 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~8 .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [1]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [3]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0 .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0 .mask = 16'h0001;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [4]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [6]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [5]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1 .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1 .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1 .mask = 16'h0001;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2 (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2 .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2 .mask = 16'hF000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [0]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [1]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [1]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~0 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~0 .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~0 .mask = 16'h1428;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~1 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [3]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [2]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [2]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~1_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~1 .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~1 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~1 .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~1 .mask = 16'h1428;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~1 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~1 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~1 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~1 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~1 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~2 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [5]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [4]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [4]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~2_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~2 .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~2 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~2 .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~2 .mask = 16'h1428;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~2 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~2 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~2 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~2 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~2 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~3 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [7]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [6]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [7]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~3_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~3 .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~3 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~3 .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~3 .mask = 16'h1248;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~3 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~3 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~3 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~3 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~3 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~1_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~2_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~3_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4 .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4 .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4 .mask = 16'h8000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|base_address~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0] .mask = 16'h0FF0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|collecting_post_data_var~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var .mask = 16'h0015;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~q ),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done .mask = 16'hFCF0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~1_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~1_combout ),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~2_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped .mask = 16'h00F4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:is_buffer_wrapped .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~0_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0] .mask = 16'h000C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~2_combout ),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1] .mask = 16'h000A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~4_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0_combout ),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~2_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2] .mask = 16'h0022;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~6_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~3_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3] .mask = 16'h0030;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~8_combout ),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~4_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4] .mask = 16'h000A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~10_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~5_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5] .mask = 16'h0300;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~12_combout ),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~6_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6] .mask = 16'h000A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~0_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(SyncReset_X16_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y14_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~0_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~1 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0] .mask = 16'h33CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[0] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~1_combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~1 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(SyncReset_X16_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y14_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~2_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~3 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1] .mask = 16'h3C3F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[1] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~2_combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~3 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(SyncReset_X16_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y14_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~4_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~5 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2] .mask = 16'hC30C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[2] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~3_combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~5 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(SyncReset_X16_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y14_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~6_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~7 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3] .mask = 16'h3C3F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[3] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~4_combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~7 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(SyncReset_X16_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y14_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~8_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~9 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4] .mask = 16'hC30C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[4] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~5_combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~9 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(SyncReset_X16_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y14_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~10_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~11 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5] .mask = 16'h3C3F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[5] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~6_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6]~q ),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~11 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X16_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y14_SIG ),
	.SyncReset(SyncReset_X16_Y14_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y14_VCC),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~12_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6] .mask = 16'hF00F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:next_address[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var .mask = 16'hCDCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[0] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter~6_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [0]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X23_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter~5_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[0] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[0] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[0] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[0] .mask = 16'hFCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[1] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~2_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [1]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~4_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[1] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[1] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[1] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[1] .mask = 16'hC0C0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~5_combout ),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [2]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X23_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~7_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[2] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[2] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[2] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[2] .mask = 16'hAA00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~8_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [3]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X23_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~10_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3] .mask = 16'hF000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4 .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4 .mask = 16'h440B;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[4] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~11_combout ),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [4]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X23_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~13_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[4] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[4] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[4] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[4] .mask = 16'hAA00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[5] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~14_combout ),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [5]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X23_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~16_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[5] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[5] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[5] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[5] .mask = 16'hAA00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[6] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~17_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [6]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X23_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~19_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[6] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[6] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[6] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[6] .mask = 16'hF000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[7] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~20_combout ),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[3]~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [7]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X23_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X23_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add3~22_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter [7]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[7] .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[7] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[7] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[7] .mask = 16'hCC00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|counter[7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~1 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~q ),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~1_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~1 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~1 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~1 .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~1 .mask = 16'hAA00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~1 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~1 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~1 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~1 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~1 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|trigger_config_deserialize|dffs [0]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|builtin:ela_trigger_flow_mgr_entity|last_level_delayed~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4 .coord_x = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4 .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4 .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4 .mask = 16'h5400;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:base_address[0]~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0_combout ),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~q ),
	.Clk(\clk~inputclkctrl_outclk_X21_Y18_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig .mask = 16'hF9F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|done~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~0 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~0 .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~0 .mask = 16'h0A08;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~4_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~0_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~6_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~0 .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~0 .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~0 .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~0 .mask = 16'h8000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~1 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~12_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~10_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Add2~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~1_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~1 .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~1 .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~1 .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~1 .mask = 16'h8000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~1 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~1 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~1 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~1 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped~1 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [0]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0_combout_X17_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|condition_delay_reg [3]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0 .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0 .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0 .mask = 16'h0088;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[1] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~1_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [1]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0_combout_X17_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[1] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[1] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[1] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[2] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~2_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [2]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0_combout_X17_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[2]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[2] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[2] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[2] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[2] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[3] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~3_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [3]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0_combout_X17_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[3]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[3] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[3] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[3] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[3] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~4_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [4]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0_combout_X17_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[4]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[4] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[4] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[4] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~5_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [5]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0_combout_X17_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[5]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[5] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[5] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[5] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[5] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[6] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|offset_count~6_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [6]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0_combout_X17_Y14_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[6]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[6] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[6] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[6] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [0]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [0]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X22_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X22_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[0]~21_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[0] .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[0] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[0] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[0] .mask = 16'h00FF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [1]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [1]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X24_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1]~7_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1]~8 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1] .mask = 16'h9911;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [2]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[1]~8 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [2]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X24_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2]~9_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2]~10 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2] .mask = 16'h5AAF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[2]~10 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [3]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X24_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3]~11_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3]~12 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3] .mask = 16'hA505;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[3]~12 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [4]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X24_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4]~13_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4]~14 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4] .mask = 16'hC33F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[4]~14 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [5]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X24_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5]~15_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5]~16 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5] .mask = 16'hC303;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_offset_config_deserialize|dffs [6]),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[5]~16 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [6]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X24_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6]~17_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6]~18 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6] .mask = 16'h3CCF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[6]~18 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [7]),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X24_Y19_SIG_SIG ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X24_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[7]~19_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count [7]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[7] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[7] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[7] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[7] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[7] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|modified_post_count[7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal1~4_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0 .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0 .mask = 16'h5054;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|process_0~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~1_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|Equal0~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0 .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0 .mask = 16'h1500;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|segment_shift_var~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~q ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on~combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on .mask = 16'hF0D0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~1 (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed~q ),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:done~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~1_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~1 .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~1 .coord_y = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~1 .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~1 .mask = 16'hCCFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~1 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~1 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~1 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~1 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~1 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [1]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on~combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:collecting_post_data_var~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[0] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[0] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[0] .mask = 16'hAC0C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[10] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [11]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [10]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~11_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [10]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[10] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[10] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[10] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[10] .mask = 16'h04CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[10] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[10] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[10] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[10] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[10] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[11] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [12]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [11]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~12_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [11]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[11] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[11] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[11] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[11] .mask = 16'h222A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[11] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[11] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[11] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[11] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[11] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[12] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [13]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [12]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~13_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [12]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[12] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[12] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[12] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[12] .mask = 16'h04CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[12] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[12] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[12] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[12] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[12] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[13] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [14]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [13]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~14_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [13]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[13] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[13] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[13] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[13] .mask = 16'h222A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[13] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[13] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[13] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[13] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[13] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[14] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [15]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [14]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~15_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [14]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[14] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[14] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[14] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[14] .mask = 16'h04CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[14] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[14] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[14] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[14] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[14] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[15] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [16]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [15]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~16_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [15]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[15] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[15] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[15] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[15] .mask = 16'h222A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[15] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[15] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[15] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[15] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[15] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[16] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.C(\altera_internal_jtag~TDIUTAP ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [16]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~17_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [16]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[16] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[16] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[16] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[16] .mask = 16'h10F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[16] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[16] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[16] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[16] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[16] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on~combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [2]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~1_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~2_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[1] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[1] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[1] .mask = 16'hB830;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[2] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on~combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [3]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~3_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[2] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[2] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[2] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[2] .mask = 16'hF3C0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[3] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [4]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X18_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~4_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[3] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[3] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[3] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[3] .mask = 16'h0FCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[4] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [5]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed [0]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_load_on~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~5_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[4] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[4] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[4] .mask = 16'hF0AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[5] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [6]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~6_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[5] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[5] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[5] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[5] .mask = 16'h04CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[6] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [7]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~7_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[6] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[6] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[6] .mask = 16'h04CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[7] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [8]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [7]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~8_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [7]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[7] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[7] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[7] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[7] .mask = 16'h222A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[8] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [9]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [8]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~9_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [8]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[8] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[8] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[8] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[8] .mask = 16'h04CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[8] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[8] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[8] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[8] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[8] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[9] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_3~0_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [10]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [9]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|_~10_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [9]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[9] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[9] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[9] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[9] .mask = 16'h04CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[9] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[9] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[9] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[9] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs[9] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0 .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0 .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0 .mask = 16'h5040;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~q ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0_combout ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][6]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1 .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1 .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1 .mask = 16'hF0D0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [1]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [0]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0 .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0 .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0 .mask = 16'h4000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [1]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [0]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0 .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0 .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0 .mask = 16'h0800;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset .mask = 16'hFFF7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~0 (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~0 .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~0 .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~0 .mask = 16'h000C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [0]),
	.B(vcc),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y18_GND),
	.SyncReset(SyncReset_X18_Y18_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena~combout__SyncLoad_X18_Y18_INV ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_comb_bita0~combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_comb_bita0~COUT ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[0] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[0] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[0] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[0] .mask = 16'h55AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[0] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[0] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[0] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[1] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [1]),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_comb_bita0~COUT ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y18_GND),
	.SyncReset(SyncReset_X18_Y18_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena~combout__SyncLoad_X18_Y18_INV ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_comb_bita1~combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_comb_bita1~COUT ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[1] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[1] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[1] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[1] .mask = 16'h3C3F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[1] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[1] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[1] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [2]),
	.B(vcc),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_comb_bita1~COUT ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y18_GND),
	.SyncReset(SyncReset_X18_Y18_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena~combout__SyncLoad_X18_Y18_INV ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_comb_bita2~combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[2] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[2] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[2] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[2] .mask = 16'hA5A5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[2] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[2] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|is_buffer_wrapped_once_sig~q ),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [1]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y18_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[0] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[0] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[0] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[0] .mask = 16'hAAF0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[10] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[2]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [11]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [10]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y14_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~10_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [10]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[10] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[10] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[10] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[10] .mask = 16'hCFC0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[10] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[10] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[10] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[10] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[10] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[11] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [12]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[3]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [11]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~11_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [11]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[11] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[11] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[11] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[11] .mask = 16'hE4E4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[11] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[11] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[11] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[11] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[11] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[12] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [13]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[4]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [12]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~12_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [12]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[12] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[12] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[12] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[12] .mask = 16'hE2E2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[12] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[12] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[12] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[12] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[12] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[13] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [14]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[5]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [13]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~13_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [13]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[13] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[13] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[13] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[13] .mask = 16'hFC0C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[13] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[13] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[13] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[13] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[13] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[14] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [0]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[6]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [14]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~14_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [14]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[14] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[14] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[14] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[14] .mask = 16'hFA0A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[14] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[14] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[14] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[14] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[14] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [0]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [2]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y18_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X21_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[1] .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[1] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[1] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[1] .mask = 16'hAAF0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [3]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [1]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y14_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~2_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[2] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[2] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[2] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[2] .mask = 16'hCACA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [4]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [2]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y14_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~3_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[3] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[3] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[3] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[3] .mask = 16'hCACA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[4] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [3]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [5]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y14_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~4_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[4] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[4] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[4] .mask = 16'hACAC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[5] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [6]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [4]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y14_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~5_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[5] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[5] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[5] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[5] .mask = 16'hCACA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[6] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [5]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [7]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y14_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~6_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[6] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[6] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[6] .mask = 16'hACAC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[7] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig [6]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [8]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [7]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y14_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~7_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [7]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[7] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[7] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[7] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[7] .mask = 16'hACAC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[8] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [9]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[0]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [8]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y14_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~8_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [8]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[8] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[8] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[8] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[8] .mask = 16'hFA0A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[8] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[8] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[8] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[8] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[8] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[9] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [10]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:last_trigger_address_var[1]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [9]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y14_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|_~9_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [9]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[9] .coord_x = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[9] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[9] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[9] .mask = 16'hFA0A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[9] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[9] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[9] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[9] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs[9] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena~combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena .mask = 16'h2000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [1]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [0]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[0] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[0] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[0] .mask = 16'hF0AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [1]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [2]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[1] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[1] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[1] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [3]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [2]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~2_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[2] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[2] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[2] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[2] .mask = 16'hCCAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [4]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [3]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~3_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[3] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[3] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[3] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[3] .mask = 16'hF0AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[4] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [5]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [4]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~4_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[4] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[4] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[4] .mask = 16'hF0CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[5] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [6]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [5]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~5_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[5] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[5] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[5] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[5] .mask = 16'hF0AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[6] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [7]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [6]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~6_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[6] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[6] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[6] .mask = 16'hF0AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[7] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [7]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [7]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X16_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|_~7_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs [7]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[7] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[7] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[7] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[7] .mask = 16'hF0FF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_data_shift_out|dffs[7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [0]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [1]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena~combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load~combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load .mask = 16'h8F0F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|ram_shift_load .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [0]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [1]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|adv_point_3_and_more:advance_pointer_counter|auto_generated|counter_reg_bit [2]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena~combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena .mask = 16'hFF40;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [0]),
	.B(vcc),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena~combout_X16_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y17_GND),
	.SyncReset(SyncReset_X16_Y17_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~combout__SyncLoad_X16_Y17_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita0~combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita0~COUT ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[0] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[0] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[0] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[0] .mask = 16'h55AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[0] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[0] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[0] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[1] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [1]),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita0~COUT ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena~combout_X16_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y17_GND),
	.SyncReset(SyncReset_X16_Y17_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~combout__SyncLoad_X16_Y17_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita1~combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita1~COUT ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[1] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[1] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[1] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[1] .mask = 16'h3C3F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[1] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[1] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[1] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[2] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [2]),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita1~COUT ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena~combout_X16_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y17_GND),
	.SyncReset(SyncReset_X16_Y17_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~combout__SyncLoad_X16_Y17_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita2~combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita2~COUT ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[2] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[2] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[2] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[2] .mask = 16'hC30C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[2] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[2] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[2] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[3] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [3]),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita2~COUT ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena~combout_X16_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y17_GND),
	.SyncReset(SyncReset_X16_Y17_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~combout__SyncLoad_X16_Y17_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita3~combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita3~COUT ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[3] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[3] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[3] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[3] .mask = 16'h3C3F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[3] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[3] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[3] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[4] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [4]),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita3~COUT ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena~combout_X16_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y17_GND),
	.SyncReset(SyncReset_X16_Y17_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~combout__SyncLoad_X16_Y17_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita4~combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita4~COUT ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[4] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[4] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[4] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[4] .mask = 16'hC30C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[4] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[4] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[4] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[5] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [5]),
	.B(vcc),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita4~COUT ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena~combout_X16_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y17_GND),
	.SyncReset(SyncReset_X16_Y17_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~combout__SyncLoad_X16_Y17_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita5~combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita5~COUT ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[5] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[5] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[5] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[5] .mask = 16'h5A5F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[5] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[5] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[5] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[6] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [6]),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita5~COUT ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena~combout_X16_Y17_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y17_GND),
	.SyncReset(SyncReset_X16_Y17_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~combout__SyncLoad_X16_Y17_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_comb_bita6~combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[6] .coord_x = 17;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[6] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[6] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[6] .mask = 16'hC3C3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[6] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[6] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~0 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~COUT ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~0 .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~0 .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~0 .mask = 16'h0F0F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~0 .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[0] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [0]),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y20_SIG_VCC ),
	.AsyncReset(AsyncReset_X17_Y20_GND),
	.SyncReset(SyncReset_X17_Y20_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0_combout__SyncLoad_X17_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita0~combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita0~COUT ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[0] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[0] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[0] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[0] .mask = 16'h33CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[0] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[0] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[0] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[1] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [1]),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita0~COUT ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y20_SIG_VCC ),
	.AsyncReset(AsyncReset_X17_Y20_GND),
	.SyncReset(SyncReset_X17_Y20_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0_combout__SyncLoad_X17_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita1~combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita1~COUT ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[1] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[1] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[1] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[1] .mask = 16'h3C3F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[1] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[1] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[1] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [2]),
	.B(vcc),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita1~COUT ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y20_SIG_VCC ),
	.AsyncReset(AsyncReset_X17_Y20_GND),
	.SyncReset(SyncReset_X17_Y20_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0_combout__SyncLoad_X17_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita2~combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita2~COUT ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[2] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[2] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[2] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[2] .mask = 16'hA50A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[2] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[2] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[2] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [3]),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita2~COUT ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y20_SIG_VCC ),
	.AsyncReset(AsyncReset_X17_Y20_GND),
	.SyncReset(SyncReset_X17_Y20_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0_combout__SyncLoad_X17_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~COUT ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3] .mask = 16'h3C3F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_comb_bita3~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0 .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0 .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0 .mask = 16'hFFFD;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [1]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [0]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y19_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[0] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[0] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[0] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[0] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[10] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [10]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [11]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [10]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y18_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~10_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [10]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[10] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[10] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[10] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[10] .mask = 16'hCCAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[10] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[10] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[10] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[10] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[10] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[11] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [12]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [11]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [11]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y18_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~11_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [11]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[11] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[11] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[11] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[11] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[11] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[11] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[11] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[11] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[11] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[12] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [13]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [12]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [12]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y18_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~12_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [12]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[12] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[12] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[12] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[12] .mask = 16'hAAF0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[12] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[12] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[12] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[12] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[12] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[13] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [13]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [14]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [13]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y18_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~13_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [13]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[13] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[13] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[13] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[13] .mask = 16'hCCAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[13] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[13] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[13] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[13] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[13] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[14] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [14]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [14]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y18_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~14_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [14]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[14] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[14] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[14] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[14] .mask = 16'hAABA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[14] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[14] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[14] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[14] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[14] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [1]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y19_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[1] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[1] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[1] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[1] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [3]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y19_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~2_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[2] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[2] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[2] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[2] .mask = 16'hCCAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [3]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [4]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y19_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~3_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[3] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[3] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[3] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[3] .mask = 16'hCCAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[4] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [5]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [4]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y19_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~4_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[4] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[4] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[4] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[4] .mask = 16'hCCF0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[5] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [6]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [5]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y19_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~5_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[5] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[5] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[5] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[5] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[6] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [7]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [6]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y19_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~6_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[6] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[6] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[6] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[6] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[7] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [7]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [8]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [7]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y19_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y19_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~7_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [7]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[7] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[7] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[7] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[7] .mask = 16'hF0AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[8] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [9]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [8]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [8]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y18_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~8_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [8]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[8] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[8] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[8] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[8] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[8] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[8] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[8] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[8] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[8] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[9] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [10]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [9]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [9]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y18_SIG_VCC ),
	.AsyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|reset_all~clkctrl_outclk__AsyncReset_X17_Y18_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|_~9_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs [9]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[9] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[9] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[9] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[9] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[9] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[9] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[9] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[9] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_data_shift_out|dffs[9] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal3~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0 .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0 .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0 .mask = 16'h000A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_ram_shift_load~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~0 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~COUT ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~0 .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~0 .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~0 .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~0 .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit [0]),
	.C(\auto_signaltap_0|~GND~combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0_combout_X18_Y20_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y20_GND),
	.SyncReset(SyncReset_X18_Y20_GND),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0_combout__SyncLoad_X18_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~COUT ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0] .mask = 16'h33CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~0_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit [0]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_comb_bita0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0 .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0 .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0 .mask = 16'hFF7F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(SyncReset_X16_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y19_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [2]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(SyncReset_X16_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y18_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [3]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(SyncReset_X16_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y18_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [4]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [5]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(SyncReset_X16_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y18_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [6]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [0]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [1]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(SyncReset_X16_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y19_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [2]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [3]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [4]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [5]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [6]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [0]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [1]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|segment_wrapped_delayed~q ),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(SyncReset_X16_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y19_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [2]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(SyncReset_X16_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y18_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [3]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(SyncReset_X16_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y18_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [4]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [5]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(SyncReset_X16_Y18_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y18_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [6]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [0]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2] (
	.A(),
	.B(),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [1]),
	.D(),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(SyncReset_X16_Y19_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y19_VCC),
	.LutOut(),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2] .mask = 16'hFFFF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [2]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [3]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [4]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [5]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|last_trigger_address_delayed [6]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [0]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8] .mask = 16'hFF00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [1]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9]~q ),
	.Clk(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X16_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9]~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9] .coord_x = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9] .mask = 16'hF0F0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|current_segment_delayed [0]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|buffer_manager:segment_shift_var~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0 .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0 .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0 .mask = 16'hA080;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][0]~q ),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][0]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[0]~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[0] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[0] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[0] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[0] .mask = 16'hFA0A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[10] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][10]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][10]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [10]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[10]~10_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [10]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[10] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[10] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[10] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[10] .mask = 16'hF0CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[10] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[10] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[10] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[10] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[10] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[11] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][11]~q ),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][11]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [11]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[11]~11_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [11]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[11] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[11] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[11] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[11] .mask = 16'hF0AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[11] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[11] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[11] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[11] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[11] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[12] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][12]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][12]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [12]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[12]~12_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [12]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[12] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[12] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[12] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[12] .mask = 16'hCCF0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[12] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[12] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[12] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[12] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[12] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[13] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][13]~q ),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][13]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [13]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[13]~13_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [13]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[13] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[13] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[13] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[13] .mask = 16'hF0AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[13] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[13] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[13] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[13] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[13] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[14] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][14]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][14]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [14]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[14]~14_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [14]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[14] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[14] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[14] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[14] .mask = 16'hF0CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[14] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[14] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[14] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[14] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[14] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][1]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][1]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[1]~1_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[1] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[1] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[1] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[1] .mask = 16'hFA50;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][2]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][2]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[2]~2_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[2] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[2] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[2] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[2] .mask = 16'hF5A0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[3] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][3]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][3]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[3]~3_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[3] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[3] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[3] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[3] .mask = 16'hFC0C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[4] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][4]~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][4]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[4]~4_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[4] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[4] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[4] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[4] .mask = 16'hCACA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[5] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][5]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][5]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[5]~5_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[5] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[5] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[5] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[5] .mask = 16'hFC0C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[6] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][6]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][6]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[6]~6_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[6] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[6] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[6] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[6] .mask = 16'hF5A0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[7] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][7]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][7]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [7]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y19_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[7]~7_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [7]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[7] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[7] .coord_y = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[7] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[7] .mask = 16'hFC0C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[8] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][8]~q ),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][8]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [8]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[8]~8_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [8]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[8] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[8] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[8] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[8] .mask = 16'hF0AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[8] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[8] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[8] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[8] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[8] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[9] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[0][9]~q ),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|cells[1][9]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [9]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X17_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|mux|auto_generated|result_node[9]~9_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq [9]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[9] .coord_x = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[9] .coord_y = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[9] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[9] .mask = 16'hF0AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[9] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[9] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[9] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[9] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xq[9] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr[0] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X18_Y20_SIG_SIG ),
	.AsyncReset(AsyncReset_X18_Y20_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr[0]~feeder_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr[0] .coord_x = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr[0] .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr[0] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr[0] .mask = 16'hCCCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|xraddr[0] .CarryEnb = 1'b1;

alta_bram9k \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 (
	.DataInA({vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc, \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][7]~q , \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][6]~q , \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][5]~q , \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][4]~q , \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][3]~q , \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][2]~q , \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][1]~q , \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|acq_data_in_pipe_reg[3][0]~q }),
	.DataInB({vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc, vcc}),
	.AddressA({\auto_hub|~GND~combout , \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [6], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [5], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [4], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [3], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [2], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [1], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_address_delayed [0], vcc, vcc, vcc, vcc, vcc}),
	.AddressB({\auto_hub|~GND~combout , \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [6], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [5], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [4], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [3], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [2], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [1], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter|auto_generated|counter_reg_bit [0], vcc, vcc, vcc, vcc, vcc}),
	.ByteEnA({vcc, vcc}),
	.ByteEnB({vcc, vcc}),
	.DataOutA({\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [17], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [16], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [15], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [14], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [13], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [12], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [11], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [10], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [9], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [8], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [7], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [6], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [5], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [4], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [3], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [2], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [1], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutA [0]}),
	.DataOutB({\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [17], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [16], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [15], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [14], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [13], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [12], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [11], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [10], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [9], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [8], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [7], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [6], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [5], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [4], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [3], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [2], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [1], \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0__DataOutB [0]}),
	.Clk0(\clk~inputclkctrl_outclk ),
	.ClkEn0(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed~q ),
	.AsyncReset0(gnd),
	.Clk1(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.AsyncReset1(gnd),
	.WeA(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|buffer_write_enable_delayed~q ),
	.ReA(gnd),
	.WeB(gnd),
	.ReB(vcc),
	.AddressStallA(gnd),
	.AddressStallB(gnd));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .coord_x = 18;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .CLKMODE = 2'b10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PACKEDMODE = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTA_CLKIN_EN = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTA_CLKOUT_EN = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTB_CLKIN_EN = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTB_CLKOUT_EN = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTA_RSTIN_EN = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTA_RSTOUT_EN = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTB_RSTIN_EN = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTB_RSTOUT_EN = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTA_WIDTH = 5'b10000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTB_WIDTH = 5'b10000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTA_WRITETHRU = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTB_WRITETHRU = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTA_OUTREG = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .PORTB_OUTREG = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .RSEN_DLY = 2'b00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .DLYTIME = 2'b00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:stp_buffer_ram|auto_generated|ram_block1a0 .INIT_VAL = 9216'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [1]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X22_Y18_SIG_INV ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[0] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[0] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[0] .mask = 16'h2112;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[0] .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[10] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [11]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [10]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X19_Y18_SIG_INV ),
	.AsyncReset(AsyncReset_X19_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~11_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [10]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[10] .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[10] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[10] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[10] .mask = 16'h0A0A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[10] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[10] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[10] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[10] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[10] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[11] (
	.A(vcc),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [12]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [11]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X19_Y18_SIG_INV ),
	.AsyncReset(AsyncReset_X19_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~12_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [11]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[11] .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[11] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[11] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[11] .mask = 16'h0F00;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[11] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[11] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[11] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[11] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[11] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [0]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [12]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X22_Y18_SIG_INV ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~13_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [12]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12] .mask = 16'h0066;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1 .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1 .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1 .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1 .mask = 16'h5540;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [2]),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X22_Y18_SIG_INV ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~2_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[1] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[1] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[1] .mask = 16'h00AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[2] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [3]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X22_Y18_SIG_INV ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~3_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[2] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[2] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[2] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[2] .mask = 16'h00CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [4]),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X22_Y18_SIG_INV ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~4_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[3] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[3] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[3] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[3] .mask = 16'h00AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[4] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [5]),
	.B(vcc),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X22_Y18_SIG_INV ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~5_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[4] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[4] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[4] .mask = 16'h00AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[5] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [6]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [0]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X22_Y18_SIG_INV ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~6_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[5] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[5] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[5] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[5] .mask = 16'h0096;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[6] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [7]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X22_Y18_SIG_INV ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~7_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[6] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[6] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[6] .mask = 16'h3300;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[7] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [8]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [7]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X19_Y18_SIG_INV ),
	.AsyncReset(AsyncReset_X19_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~8_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [7]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[7] .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[7] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[7] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[7] .mask = 16'h4444;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[8] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [9]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [8]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X19_Y18_SIG_INV ),
	.AsyncReset(AsyncReset_X19_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~9_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [8]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[8] .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[8] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[8] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[8] .mask = 16'h0A0A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[8] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[8] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[8] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[8] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[8] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[9] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [10]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [9]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X19_Y18_SIG_INV ),
	.AsyncReset(AsyncReset_X19_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr~10_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [9]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[9] .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[9] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[9] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[9] .mask = 16'h0A0A;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[9] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[9] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[9] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[9] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[9] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9]~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0 .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0 .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0 .mask = 16'h0200;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen~0 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [0]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [1]),
	.D(vcc),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0]~32_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0]~33 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0] .mask = 16'h55AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [10]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [11]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9]~53 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [10]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~54_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~55 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [10]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10] .mask = 16'h3CCF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~34 (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8]~q ),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~34_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~34 .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~34 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~34 .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~34 .mask = 16'h3F3F;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~34 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~34 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~34 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~34 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~34 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~34_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sdr~combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~9_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|LessThan0~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35 .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35 .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35 .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35 .mask = 16'hA888;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [11]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [12]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~55 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [11]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11]~56_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11]~57 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [11]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11] .mask = 16'hA505;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [12]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [13]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[11]~57 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [12]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12]~58_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12]~59 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [12]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12] .mask = 16'h5AAF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [13]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [14]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[12]~59 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [13]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13]~60_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13]~61 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [13]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13] .mask = 16'hA505;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [14]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [15]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[13]~61 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [14]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14]~62_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14]~63 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [14]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14] .mask = 16'h3CCF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [15]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [16]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[14]~63 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [15]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15]~64_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15]~65 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [15]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15] .mask = 16'hC303;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [16]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [17]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[15]~65 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [16]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16]~66_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16]~67 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [16]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16] .mask = 16'h5AAF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [17]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [18]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[16]~67 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [17]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17]~68_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17]~69 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [17]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17] .mask = 16'hC303;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [18]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [19]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[17]~69 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [18]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18]~70_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18]~71 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [18]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18] .mask = 16'h3CCF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [19]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [20]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[18]~71 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [19]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19]~72_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19]~73 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [19]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19] .mask = 16'hA505;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [1]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [2]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[0]~33 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1]~36_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1]~37 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1] .mask = 16'hC303;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [20]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [21]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[19]~73 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [20]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20]~74_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20]~75 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [20]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20] .mask = 16'h5AAF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [21]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [22]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[20]~75 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [21]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21]~76_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21]~77 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [21]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21] .mask = 16'hA505;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [22]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [23]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[21]~77 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [22]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22]~78_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22]~79 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [22]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22] .mask = 16'h5AAF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [23]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [24]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[22]~79 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [23]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23]~80_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23]~81 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [23]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23] .mask = 16'hC303;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [24]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [25]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[23]~81 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [24]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24]~82_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24]~83 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [24]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24] .mask = 16'h3CCF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [25]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [26]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[24]~83 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [25]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25]~84_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25]~85 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [25]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25] .mask = 16'hC303;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [26]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [27]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[25]~85 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [26]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26]~86_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26]~87 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [26]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26] .mask = 16'h5AAF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [27]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [28]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[26]~87 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [27]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27]~88_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27]~89 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [27]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27] .coord_z = 11;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27] .mask = 16'hC303;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [28]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [29]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[27]~89 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [28]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28]~90_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28]~91 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [28]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28] .mask = 16'h3CCF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [29]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [30]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[28]~91 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [29]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29]~92_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29]~93 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [29]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29] .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29] .mask = 16'hA505;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [2]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [3]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[1]~37 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2]~38_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2]~39 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2] .mask = 16'h3CCF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [30]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [31]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[29]~93 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [30]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30]~94_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30]~95 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [30]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30] .mask = 16'h5AAF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[31] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [31]),
	.B(vcc),
	.C(\altera_internal_jtag~TDIUTAP ),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[30]~95 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [31]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y19_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[31]~96_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [31]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[31] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[31] .coord_y = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[31] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[31] .mask = 16'hA5A5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[31] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[31] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[31] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[31] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[31] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [3]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [4]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[2]~39 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3]~40_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3]~41 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3] .coord_z = 3;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3] .mask = 16'hA505;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [4]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [5]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[3]~41 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4]~42_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4]~43 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4] .mask = 16'h5AAF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [5]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [6]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[4]~43 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5]~44_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5]~45 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5] .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5] .mask = 16'hA505;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [6]),
	.B(vcc),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [7]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[5]~45 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6]~46_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6]~47 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6] .mask = 16'h5AAF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [7]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [8]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[6]~47 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [7]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7]~48_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7]~49 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [7]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7] .mask = 16'hC303;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [8]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [9]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[7]~49 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [8]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8]~50_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8]~51 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [8]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8] .mask = 16'h3CCF;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [9]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [10]),
	.D(vcc),
	.Cin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[8]~51 ),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [9]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ),
	.AsyncReset(AsyncReset_X14_Y20_GND),
	.SyncReset(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ),
	.ShiftData(),
	.SyncLoad(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9]~52_combout ),
	.Cout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9]~53 ),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [9]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9] .coord_y = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9] .mask = 16'hC303;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9] .modeMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9] .BypassEn = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[9] .CarryEnb = 1'b0;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [1]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [0]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [0]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X22_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [0]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0] .mask = 16'hCCAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1 (
	.A(vcc),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9]~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~0_combout ),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1 .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1 .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1 .mask = 16'hC0C0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[10] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [10]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [11]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [10]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X19_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~11_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [10]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[10] .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[10] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[10] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[10] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[10] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[10] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[10] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[10] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[10] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[11] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [11]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [12]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [11]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X19_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~12_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [11]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[11] .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[11] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[11] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[11] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[11] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[11] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[11] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[11] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[11] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[12] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [13]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [12]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [12]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X19_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~13_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [12]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[12] .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[12] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[12] .coord_z = 12;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[12] .mask = 16'hEE44;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[12] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[12] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[12] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[12] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[12] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[13] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [14]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [13]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X19_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~14_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [13]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[13] .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[13] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[13] .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[13] .mask = 16'hA2AA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[13] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[13] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[13] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[13] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[13] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[14] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [15]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [14]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X19_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~15_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [14]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[14] .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[14] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[14] .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[14] .mask = 16'h8CCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[14] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[14] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[14] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[14] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[14] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[15] (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.B(\altera_internal_jtag~TDIUTAP ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [15]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X19_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~16_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [15]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[15] .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[15] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[15] .coord_z = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[15] .mask = 16'h8CCC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[15] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[15] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[15] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[15] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[15] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[1] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [1]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [2]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [1]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X22_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~2_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [1]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[1] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[1] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[1] .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[1] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[1] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[1] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[1] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[1] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[1] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[2] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [2]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [3]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [2]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X22_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~3_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [2]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[2] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[2] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[2] .coord_z = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[2] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[2] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[2] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[2] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[2] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[2] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[3] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [4]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [3]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [3]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X22_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~4_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [3]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[3] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[3] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[3] .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[3] .mask = 16'hCCAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[3] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[3] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[3] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[3] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[3] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[4] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [4]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [5]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [4]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X22_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~5_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [4]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[4] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[4] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[4] .coord_z = 0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[4] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[4] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[4] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[4] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[4] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[4] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[5] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [5]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [6]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [5]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X22_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~6_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [5]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[5] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[5] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[5] .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[5] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[5] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[5] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[5] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[5] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[5] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[6] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [6]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [7]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [6]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X22_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~7_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [6]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[6] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[6] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[6] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[6] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[6] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[6] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[6] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[6] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[6] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[7] (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [7]),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [8]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [7]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X22_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~8_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [7]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[7] .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[7] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[7] .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[7] .mask = 16'hCCF0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[7] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[7] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[7] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[7] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[7] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[8] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [9]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [8]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [8]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X19_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~9_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [8]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[8] .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[8] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[8] .coord_z = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[8] .mask = 16'hCCAA;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[8] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[8] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[8] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[8] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[8] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[9] (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr [9]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [10]),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|cdr~0_combout ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [9]),
	.Clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X19_Y18_SIG_SIG ),
	.AsyncReset(AsyncReset_X19_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg~10_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [9]));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[9] .coord_x = 7;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[9] .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[9] .coord_z = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[9] .mask = 16'hAACC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[9] .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[9] .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[9] .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[9] .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[9] .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~1 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg [0]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~0_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9]~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~1_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~1 .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~1 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~1 .coord_z = 14;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~1 .mask = 16'h0A0C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~1 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~1 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~1 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~1 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~1 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2 (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][8]~q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9]~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2 .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2 .coord_z = 2;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2 .mask = 16'h0001;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~3 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|info_data_shift_out|dffs [0]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR [0]),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~3_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~3 .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~3 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~3 .coord_z = 6;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~3 .mask = 16'hACA0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~3 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~3 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~3 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~3 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~3 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~4 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg [0]),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][9]~q ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~4_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~4 .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~4 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~4 .coord_z = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~4 .mask = 16'hECA0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~4 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~4 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~4 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~4 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~4 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~5 (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|bypass_reg_out~q ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_register|dffs [0]),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~5_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~5 .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~5 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~5 .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~5 .mask = 16'hF0CC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~5 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~5 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~5 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~5 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~5 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~6 (
	.A(vcc),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~2_combout ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][5]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~6_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~6 .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~6 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~6 .coord_z = 1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~6 .mask = 16'h000C;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~6 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~6 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~6 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~6 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~6 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7 (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~5_combout ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~4_combout ),
	.C(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~6_combout ),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7_combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7 .coord_x = 9;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7 .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7 .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7 .mask = 16'hFFEC;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7 .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7 .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7 .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7 .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_internal~7 .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|run~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~2_combout ),
	.C(vcc),
	.D(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff~q ),
	.Clk(\clk~inputclkctrl_outclk_X18_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff .coord_z = 4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff .mask = 16'h75A8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_ff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff (
	.A(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|power_up_mode_source_reg~q ),
	.B(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|ela_control|trigger_config_deserialize|dffs [0]),
	.C(vcc),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.Cin(),
	.Qin(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff~q ),
	.Clk(\clk~inputclkctrl_outclk_X18_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X18_Y19_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff~0_combout ),
	.Cout(),
	.Q(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff~q ));
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff .coord_x = 10;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff .coord_y = 15;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff .coord_z = 13;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff .mask = 16'hCCE4;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff .FeedbackMux = 1'b1;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_out_mode_ff .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena (
	.A(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.B(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.C(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.D(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena .coord_x = 8;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena .coord_y = 16;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena .coord_z = 5;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena .mask = 16'h2000;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena .modeMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena .ShiftMux = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena .BypassEn = 1'b0;
defparam \auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena .CarryEnb = 1'b1;

alta_slice \auto_signaltap_0|~GND (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\auto_signaltap_0|~GND~combout ),
	.Cout(),
	.Q());
defparam \auto_signaltap_0|~GND .coord_x = 17;
defparam \auto_signaltap_0|~GND .coord_y = 16;
defparam \auto_signaltap_0|~GND .coord_z = 4;
defparam \auto_signaltap_0|~GND .mask = 16'h0000;
defparam \auto_signaltap_0|~GND .modeMux = 1'b0;
defparam \auto_signaltap_0|~GND .FeedbackMux = 1'b0;
defparam \auto_signaltap_0|~GND .ShiftMux = 1'b0;
defparam \auto_signaltap_0|~GND .BypassEn = 1'b0;
defparam \auto_signaltap_0|~GND .CarryEnb = 1'b1;

alta_dio \cam_data[0]~input (
	.padio(cam_data[0]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[0]~input_o ),
	.regout());
defparam \cam_data[0]~input .coord_x = 11;
defparam \cam_data[0]~input .coord_y = 0;
defparam \cam_data[0]~input .coord_z = 1;
defparam \cam_data[0]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[0]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[0]~input .IN_POWERUP = 1'b0;
defparam \cam_data[0]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[0]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[0]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[0]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[0]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[0]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[0]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[0]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[0]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[0]~input .OUT_DDIO = 1'b0;
defparam \cam_data[0]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[0]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[0]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[0]~input .OE_POWERUP = 1'b0;
defparam \cam_data[0]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[0]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[0]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[0]~input .OE_DDIO = 1'b0;
defparam \cam_data[0]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[0]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[0]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[0]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[0]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[0]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[0]~input .CFG_KEEP = 2'b00;
defparam \cam_data[0]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[0]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[0]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[0]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[0]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[0]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[0]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[0]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[0]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[0]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[0]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[0]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[0]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[0]~input .OUT_DELAY = 1'b0;
defparam \cam_data[0]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[0]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[1]~input (
	.padio(cam_data[1]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[1]~input_o ),
	.regout());
defparam \cam_data[1]~input .coord_x = 6;
defparam \cam_data[1]~input .coord_y = 0;
defparam \cam_data[1]~input .coord_z = 0;
defparam \cam_data[1]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[1]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[1]~input .IN_POWERUP = 1'b0;
defparam \cam_data[1]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[1]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[1]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[1]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[1]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[1]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[1]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[1]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[1]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[1]~input .OUT_DDIO = 1'b0;
defparam \cam_data[1]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[1]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[1]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[1]~input .OE_POWERUP = 1'b0;
defparam \cam_data[1]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[1]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[1]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[1]~input .OE_DDIO = 1'b0;
defparam \cam_data[1]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[1]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[1]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[1]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[1]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[1]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[1]~input .CFG_KEEP = 2'b00;
defparam \cam_data[1]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[1]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[1]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[1]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[1]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[1]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[1]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[1]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[1]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[1]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[1]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[1]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[1]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[1]~input .OUT_DELAY = 1'b0;
defparam \cam_data[1]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[1]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[2]~input (
	.padio(cam_data[2]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[2]~input_o ),
	.regout());
defparam \cam_data[2]~input .coord_x = 6;
defparam \cam_data[2]~input .coord_y = 0;
defparam \cam_data[2]~input .coord_z = 1;
defparam \cam_data[2]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[2]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[2]~input .IN_POWERUP = 1'b0;
defparam \cam_data[2]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[2]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[2]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[2]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[2]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[2]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[2]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[2]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[2]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[2]~input .OUT_DDIO = 1'b0;
defparam \cam_data[2]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[2]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[2]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[2]~input .OE_POWERUP = 1'b0;
defparam \cam_data[2]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[2]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[2]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[2]~input .OE_DDIO = 1'b0;
defparam \cam_data[2]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[2]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[2]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[2]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[2]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[2]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[2]~input .CFG_KEEP = 2'b00;
defparam \cam_data[2]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[2]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[2]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[2]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[2]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[2]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[2]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[2]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[2]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[2]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[2]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[2]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[2]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[2]~input .OUT_DELAY = 1'b0;
defparam \cam_data[2]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[2]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[3]~input (
	.padio(cam_data[3]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[3]~input_o ),
	.regout());
defparam \cam_data[3]~input .coord_x = 5;
defparam \cam_data[3]~input .coord_y = 0;
defparam \cam_data[3]~input .coord_z = 2;
defparam \cam_data[3]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[3]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[3]~input .IN_POWERUP = 1'b0;
defparam \cam_data[3]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[3]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[3]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[3]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[3]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[3]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[3]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[3]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[3]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[3]~input .OUT_DDIO = 1'b0;
defparam \cam_data[3]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[3]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[3]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[3]~input .OE_POWERUP = 1'b0;
defparam \cam_data[3]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[3]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[3]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[3]~input .OE_DDIO = 1'b0;
defparam \cam_data[3]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[3]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[3]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[3]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[3]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[3]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[3]~input .CFG_KEEP = 2'b00;
defparam \cam_data[3]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[3]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[3]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[3]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[3]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[3]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[3]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[3]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[3]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[3]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[3]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[3]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[3]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[3]~input .OUT_DELAY = 1'b0;
defparam \cam_data[3]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[3]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[4]~input (
	.padio(cam_data[4]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[4]~input_o ),
	.regout());
defparam \cam_data[4]~input .coord_x = 3;
defparam \cam_data[4]~input .coord_y = 0;
defparam \cam_data[4]~input .coord_z = 0;
defparam \cam_data[4]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[4]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[4]~input .IN_POWERUP = 1'b0;
defparam \cam_data[4]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[4]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[4]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[4]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[4]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[4]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[4]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[4]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[4]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[4]~input .OUT_DDIO = 1'b0;
defparam \cam_data[4]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[4]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[4]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[4]~input .OE_POWERUP = 1'b0;
defparam \cam_data[4]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[4]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[4]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[4]~input .OE_DDIO = 1'b0;
defparam \cam_data[4]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[4]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[4]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[4]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[4]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[4]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[4]~input .CFG_KEEP = 2'b00;
defparam \cam_data[4]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[4]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[4]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[4]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[4]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[4]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[4]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[4]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[4]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[4]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[4]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[4]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[4]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[4]~input .OUT_DELAY = 1'b0;
defparam \cam_data[4]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[4]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[5]~input (
	.padio(cam_data[5]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[5]~input_o ),
	.regout());
defparam \cam_data[5]~input .coord_x = 3;
defparam \cam_data[5]~input .coord_y = 0;
defparam \cam_data[5]~input .coord_z = 1;
defparam \cam_data[5]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[5]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[5]~input .IN_POWERUP = 1'b0;
defparam \cam_data[5]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[5]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[5]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[5]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[5]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[5]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[5]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[5]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[5]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[5]~input .OUT_DDIO = 1'b0;
defparam \cam_data[5]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[5]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[5]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[5]~input .OE_POWERUP = 1'b0;
defparam \cam_data[5]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[5]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[5]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[5]~input .OE_DDIO = 1'b0;
defparam \cam_data[5]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[5]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[5]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[5]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[5]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[5]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[5]~input .CFG_KEEP = 2'b00;
defparam \cam_data[5]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[5]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[5]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[5]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[5]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[5]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[5]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[5]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[5]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[5]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[5]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[5]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[5]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[5]~input .OUT_DELAY = 1'b0;
defparam \cam_data[5]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[5]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[6]~input (
	.padio(cam_data[6]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[6]~input_o ),
	.regout());
defparam \cam_data[6]~input .coord_x = 0;
defparam \cam_data[6]~input .coord_y = 4;
defparam \cam_data[6]~input .coord_z = 2;
defparam \cam_data[6]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[6]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[6]~input .IN_POWERUP = 1'b0;
defparam \cam_data[6]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[6]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[6]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[6]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[6]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[6]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[6]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[6]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[6]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[6]~input .OUT_DDIO = 1'b0;
defparam \cam_data[6]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[6]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[6]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[6]~input .OE_POWERUP = 1'b0;
defparam \cam_data[6]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[6]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[6]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[6]~input .OE_DDIO = 1'b0;
defparam \cam_data[6]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[6]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[6]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[6]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[6]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[6]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[6]~input .CFG_KEEP = 2'b00;
defparam \cam_data[6]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[6]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[6]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[6]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[6]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[6]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[6]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[6]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[6]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[6]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[6]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[6]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[6]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[6]~input .OUT_DELAY = 1'b0;
defparam \cam_data[6]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[6]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_data[7]~input (
	.padio(cam_data[7]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_data[7]~input_o ),
	.regout());
defparam \cam_data[7]~input .coord_x = 0;
defparam \cam_data[7]~input .coord_y = 4;
defparam \cam_data[7]~input .coord_z = 3;
defparam \cam_data[7]~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_data[7]~input .IN_SYNC_MODE = 1'b0;
defparam \cam_data[7]~input .IN_POWERUP = 1'b0;
defparam \cam_data[7]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_data[7]~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_data[7]~input .OUT_REG_MODE = 1'b0;
defparam \cam_data[7]~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_data[7]~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_data[7]~input .OUT_POWERUP = 1'b0;
defparam \cam_data[7]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_data[7]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_data[7]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_data[7]~input .OUT_DDIO = 1'b0;
defparam \cam_data[7]~input .OE_REG_MODE = 1'b0;
defparam \cam_data[7]~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_data[7]~input .OE_SYNC_MODE = 1'b0;
defparam \cam_data[7]~input .OE_POWERUP = 1'b0;
defparam \cam_data[7]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_data[7]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_data[7]~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_data[7]~input .OE_DDIO = 1'b0;
defparam \cam_data[7]~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_data[7]~input .CFG_PULL_UP = 1'b0;
defparam \cam_data[7]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_data[7]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_data[7]~input .CFG_PDRV = 7'b0011010;
defparam \cam_data[7]~input .CFG_NDRV = 7'b0011000;
defparam \cam_data[7]~input .CFG_KEEP = 2'b00;
defparam \cam_data[7]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_data[7]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_data[7]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_data[7]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_data[7]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_data[7]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_data[7]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_data[7]~input .CFG_OSCDIV = 2'b00;
defparam \cam_data[7]~input .CFG_ROCTUSR = 1'b0;
defparam \cam_data[7]~input .CFG_SEL_CUA = 1'b0;
defparam \cam_data[7]~input .CFG_ROCT_EN = 1'b0;
defparam \cam_data[7]~input .INPUT_ONLY = 1'b0;
defparam \cam_data[7]~input .DPCLK_DELAY = 4'b0000;
defparam \cam_data[7]~input .OUT_DELAY = 1'b0;
defparam \cam_data[7]~input .IN_DATA_DELAY = 3'b000;
defparam \cam_data[7]~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_hsync~input (
	.padio(cam_hsync),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_hsync~input_o ),
	.regout());
defparam \cam_hsync~input .coord_x = 0;
defparam \cam_hsync~input .coord_y = 8;
defparam \cam_hsync~input .coord_z = 2;
defparam \cam_hsync~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_hsync~input .IN_SYNC_MODE = 1'b0;
defparam \cam_hsync~input .IN_POWERUP = 1'b0;
defparam \cam_hsync~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_hsync~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_hsync~input .OUT_REG_MODE = 1'b0;
defparam \cam_hsync~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_hsync~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_hsync~input .OUT_POWERUP = 1'b0;
defparam \cam_hsync~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_hsync~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_hsync~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_hsync~input .OUT_DDIO = 1'b0;
defparam \cam_hsync~input .OE_REG_MODE = 1'b0;
defparam \cam_hsync~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_hsync~input .OE_SYNC_MODE = 1'b0;
defparam \cam_hsync~input .OE_POWERUP = 1'b0;
defparam \cam_hsync~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_hsync~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_hsync~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_hsync~input .OE_DDIO = 1'b0;
defparam \cam_hsync~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_hsync~input .CFG_PULL_UP = 1'b0;
defparam \cam_hsync~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_hsync~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_hsync~input .CFG_PDRV = 7'b0011010;
defparam \cam_hsync~input .CFG_NDRV = 7'b0011000;
defparam \cam_hsync~input .CFG_KEEP = 2'b00;
defparam \cam_hsync~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_hsync~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_hsync~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_hsync~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_hsync~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_hsync~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_hsync~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_hsync~input .CFG_OSCDIV = 2'b00;
defparam \cam_hsync~input .CFG_ROCTUSR = 1'b0;
defparam \cam_hsync~input .CFG_SEL_CUA = 1'b0;
defparam \cam_hsync~input .CFG_ROCT_EN = 1'b0;
defparam \cam_hsync~input .INPUT_ONLY = 1'b0;
defparam \cam_hsync~input .DPCLK_DELAY = 4'b0000;
defparam \cam_hsync~input .OUT_DELAY = 1'b0;
defparam \cam_hsync~input .IN_DATA_DELAY = 3'b000;
defparam \cam_hsync~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_pclk~input (
	.padio(cam_pclk),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_pclk~input_o ),
	.regout());
defparam \cam_pclk~input .coord_x = 0;
defparam \cam_pclk~input .coord_y = 8;
defparam \cam_pclk~input .coord_z = 1;
defparam \cam_pclk~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_pclk~input .IN_SYNC_MODE = 1'b0;
defparam \cam_pclk~input .IN_POWERUP = 1'b0;
defparam \cam_pclk~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_pclk~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_pclk~input .OUT_REG_MODE = 1'b0;
defparam \cam_pclk~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_pclk~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_pclk~input .OUT_POWERUP = 1'b0;
defparam \cam_pclk~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_pclk~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_pclk~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_pclk~input .OUT_DDIO = 1'b0;
defparam \cam_pclk~input .OE_REG_MODE = 1'b0;
defparam \cam_pclk~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_pclk~input .OE_SYNC_MODE = 1'b0;
defparam \cam_pclk~input .OE_POWERUP = 1'b0;
defparam \cam_pclk~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_pclk~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_pclk~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_pclk~input .OE_DDIO = 1'b0;
defparam \cam_pclk~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_pclk~input .CFG_PULL_UP = 1'b0;
defparam \cam_pclk~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_pclk~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_pclk~input .CFG_PDRV = 7'b0011010;
defparam \cam_pclk~input .CFG_NDRV = 7'b0011000;
defparam \cam_pclk~input .CFG_KEEP = 2'b00;
defparam \cam_pclk~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_pclk~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_pclk~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_pclk~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_pclk~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_pclk~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_pclk~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_pclk~input .CFG_OSCDIV = 2'b00;
defparam \cam_pclk~input .CFG_ROCTUSR = 1'b0;
defparam \cam_pclk~input .CFG_SEL_CUA = 1'b0;
defparam \cam_pclk~input .CFG_ROCT_EN = 1'b0;
defparam \cam_pclk~input .INPUT_ONLY = 1'b0;
defparam \cam_pclk~input .DPCLK_DELAY = 4'b0000;
defparam \cam_pclk~input .OUT_DELAY = 1'b0;
defparam \cam_pclk~input .IN_DATA_DELAY = 3'b000;
defparam \cam_pclk~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_pdown~output (
	.padio(cam_pdown),
	.datain(gnd),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \cam_pdown~output .coord_x = 22;
defparam \cam_pdown~output .coord_y = 0;
defparam \cam_pdown~output .coord_z = 0;
defparam \cam_pdown~output .IN_ASYNC_MODE = 1'b0;
defparam \cam_pdown~output .IN_SYNC_MODE = 1'b0;
defparam \cam_pdown~output .IN_POWERUP = 1'b0;
defparam \cam_pdown~output .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_pdown~output .IN_SYNC_DISABLE = 1'b0;
defparam \cam_pdown~output .OUT_REG_MODE = 1'b0;
defparam \cam_pdown~output .OUT_ASYNC_MODE = 1'b0;
defparam \cam_pdown~output .OUT_SYNC_MODE = 1'b0;
defparam \cam_pdown~output .OUT_POWERUP = 1'b0;
defparam \cam_pdown~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_pdown~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_pdown~output .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_pdown~output .OUT_DDIO = 1'b0;
defparam \cam_pdown~output .OE_REG_MODE = 1'b0;
defparam \cam_pdown~output .OE_ASYNC_MODE = 1'b0;
defparam \cam_pdown~output .OE_SYNC_MODE = 1'b0;
defparam \cam_pdown~output .OE_POWERUP = 1'b0;
defparam \cam_pdown~output .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_pdown~output .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_pdown~output .OE_SYNC_DISABLE = 1'b0;
defparam \cam_pdown~output .OE_DDIO = 1'b0;
defparam \cam_pdown~output .CFG_TRI_INPUT = 1'b0;
defparam \cam_pdown~output .CFG_PULL_UP = 1'b0;
defparam \cam_pdown~output .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_pdown~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_pdown~output .CFG_PDRV = 7'b0011010;
defparam \cam_pdown~output .CFG_NDRV = 7'b0011000;
defparam \cam_pdown~output .CFG_KEEP = 2'b00;
defparam \cam_pdown~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_pdown~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_pdown~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_pdown~output .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_pdown~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_pdown~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_pdown~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_pdown~output .CFG_OSCDIV = 2'b00;
defparam \cam_pdown~output .CFG_ROCTUSR = 1'b0;
defparam \cam_pdown~output .CFG_SEL_CUA = 1'b0;
defparam \cam_pdown~output .CFG_ROCT_EN = 1'b0;
defparam \cam_pdown~output .INPUT_ONLY = 1'b0;
defparam \cam_pdown~output .DPCLK_DELAY = 4'b0000;
defparam \cam_pdown~output .OUT_DELAY = 1'b0;
defparam \cam_pdown~output .IN_DATA_DELAY = 3'b000;
defparam \cam_pdown~output .IN_REG_DELAY = 3'b000;

alta_dio \cam_reset~output (
	.padio(cam_reset),
	.datain(!\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \cam_reset~output .coord_x = 22;
defparam \cam_reset~output .coord_y = 0;
defparam \cam_reset~output .coord_z = 1;
defparam \cam_reset~output .IN_ASYNC_MODE = 1'b0;
defparam \cam_reset~output .IN_SYNC_MODE = 1'b0;
defparam \cam_reset~output .IN_POWERUP = 1'b0;
defparam \cam_reset~output .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_reset~output .IN_SYNC_DISABLE = 1'b0;
defparam \cam_reset~output .OUT_REG_MODE = 1'b0;
defparam \cam_reset~output .OUT_ASYNC_MODE = 1'b0;
defparam \cam_reset~output .OUT_SYNC_MODE = 1'b0;
defparam \cam_reset~output .OUT_POWERUP = 1'b0;
defparam \cam_reset~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_reset~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_reset~output .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_reset~output .OUT_DDIO = 1'b0;
defparam \cam_reset~output .OE_REG_MODE = 1'b0;
defparam \cam_reset~output .OE_ASYNC_MODE = 1'b0;
defparam \cam_reset~output .OE_SYNC_MODE = 1'b0;
defparam \cam_reset~output .OE_POWERUP = 1'b0;
defparam \cam_reset~output .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_reset~output .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_reset~output .OE_SYNC_DISABLE = 1'b0;
defparam \cam_reset~output .OE_DDIO = 1'b0;
defparam \cam_reset~output .CFG_TRI_INPUT = 1'b0;
defparam \cam_reset~output .CFG_PULL_UP = 1'b0;
defparam \cam_reset~output .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_reset~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_reset~output .CFG_PDRV = 7'b0011010;
defparam \cam_reset~output .CFG_NDRV = 7'b0011000;
defparam \cam_reset~output .CFG_KEEP = 2'b00;
defparam \cam_reset~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_reset~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_reset~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_reset~output .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_reset~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_reset~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_reset~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_reset~output .CFG_OSCDIV = 2'b00;
defparam \cam_reset~output .CFG_ROCTUSR = 1'b0;
defparam \cam_reset~output .CFG_SEL_CUA = 1'b0;
defparam \cam_reset~output .CFG_ROCT_EN = 1'b0;
defparam \cam_reset~output .INPUT_ONLY = 1'b0;
defparam \cam_reset~output .DPCLK_DELAY = 4'b0000;
defparam \cam_reset~output .OUT_DELAY = 1'b0;
defparam \cam_reset~output .IN_DATA_DELAY = 3'b000;
defparam \cam_reset~output .IN_REG_DELAY = 3'b000;

alta_dio \cam_scl~output (
	.padio(cam_scl),
	.datain(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10_combout ),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \cam_scl~output .coord_x = 0;
defparam \cam_scl~output .coord_y = 13;
defparam \cam_scl~output .coord_z = 2;
defparam \cam_scl~output .IN_ASYNC_MODE = 1'b0;
defparam \cam_scl~output .IN_SYNC_MODE = 1'b0;
defparam \cam_scl~output .IN_POWERUP = 1'b0;
defparam \cam_scl~output .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_scl~output .IN_SYNC_DISABLE = 1'b0;
defparam \cam_scl~output .OUT_REG_MODE = 1'b0;
defparam \cam_scl~output .OUT_ASYNC_MODE = 1'b0;
defparam \cam_scl~output .OUT_SYNC_MODE = 1'b0;
defparam \cam_scl~output .OUT_POWERUP = 1'b0;
defparam \cam_scl~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_scl~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_scl~output .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_scl~output .OUT_DDIO = 1'b0;
defparam \cam_scl~output .OE_REG_MODE = 1'b0;
defparam \cam_scl~output .OE_ASYNC_MODE = 1'b0;
defparam \cam_scl~output .OE_SYNC_MODE = 1'b0;
defparam \cam_scl~output .OE_POWERUP = 1'b0;
defparam \cam_scl~output .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_scl~output .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_scl~output .OE_SYNC_DISABLE = 1'b0;
defparam \cam_scl~output .OE_DDIO = 1'b0;
defparam \cam_scl~output .CFG_TRI_INPUT = 1'b0;
defparam \cam_scl~output .CFG_PULL_UP = 1'b0;
defparam \cam_scl~output .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_scl~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_scl~output .CFG_PDRV = 7'b0011010;
defparam \cam_scl~output .CFG_NDRV = 7'b0011000;
defparam \cam_scl~output .CFG_KEEP = 2'b00;
defparam \cam_scl~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_scl~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_scl~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_scl~output .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_scl~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_scl~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_scl~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_scl~output .CFG_OSCDIV = 2'b00;
defparam \cam_scl~output .CFG_ROCTUSR = 1'b0;
defparam \cam_scl~output .CFG_SEL_CUA = 1'b0;
defparam \cam_scl~output .CFG_ROCT_EN = 1'b0;
defparam \cam_scl~output .INPUT_ONLY = 1'b0;
defparam \cam_scl~output .DPCLK_DELAY = 4'b0000;
defparam \cam_scl~output .OUT_DELAY = 1'b0;
defparam \cam_scl~output .IN_DATA_DELAY = 3'b000;
defparam \cam_scl~output .IN_REG_DELAY = 3'b000;

alta_dio \cam_sda~output (
	.padio(cam_sda),
	.datain(!\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.datainh(gnd),
	.oe(\camera_if_inst|u_I2C_AV_Config|u0|SDO~4_combout ),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_sda~input_o ),
	.regout());
defparam \cam_sda~output .coord_x = 0;
defparam \cam_sda~output .coord_y = 13;
defparam \cam_sda~output .coord_z = 1;
defparam \cam_sda~output .IN_ASYNC_MODE = 1'b0;
defparam \cam_sda~output .IN_SYNC_MODE = 1'b0;
defparam \cam_sda~output .IN_POWERUP = 1'b0;
defparam \cam_sda~output .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_sda~output .IN_SYNC_DISABLE = 1'b0;
defparam \cam_sda~output .OUT_REG_MODE = 1'b0;
defparam \cam_sda~output .OUT_ASYNC_MODE = 1'b0;
defparam \cam_sda~output .OUT_SYNC_MODE = 1'b0;
defparam \cam_sda~output .OUT_POWERUP = 1'b0;
defparam \cam_sda~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_sda~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_sda~output .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_sda~output .OUT_DDIO = 1'b0;
defparam \cam_sda~output .OE_REG_MODE = 1'b0;
defparam \cam_sda~output .OE_ASYNC_MODE = 1'b0;
defparam \cam_sda~output .OE_SYNC_MODE = 1'b0;
defparam \cam_sda~output .OE_POWERUP = 1'b0;
defparam \cam_sda~output .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_sda~output .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_sda~output .OE_SYNC_DISABLE = 1'b0;
defparam \cam_sda~output .OE_DDIO = 1'b0;
defparam \cam_sda~output .CFG_TRI_INPUT = 1'b0;
defparam \cam_sda~output .CFG_PULL_UP = 1'b0;
defparam \cam_sda~output .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_sda~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_sda~output .CFG_PDRV = 7'b0011010;
defparam \cam_sda~output .CFG_NDRV = 7'b0011000;
defparam \cam_sda~output .CFG_KEEP = 2'b00;
defparam \cam_sda~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_sda~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_sda~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_sda~output .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_sda~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_sda~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_sda~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_sda~output .CFG_OSCDIV = 2'b00;
defparam \cam_sda~output .CFG_ROCTUSR = 1'b0;
defparam \cam_sda~output .CFG_SEL_CUA = 1'b0;
defparam \cam_sda~output .CFG_ROCT_EN = 1'b0;
defparam \cam_sda~output .INPUT_ONLY = 1'b0;
defparam \cam_sda~output .DPCLK_DELAY = 4'b0000;
defparam \cam_sda~output .OUT_DELAY = 1'b0;
defparam \cam_sda~output .IN_DATA_DELAY = 3'b000;
defparam \cam_sda~output .IN_REG_DELAY = 3'b000;

alta_dio \cam_vsync~input (
	.padio(cam_vsync),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\cam_vsync~input_o ),
	.regout());
defparam \cam_vsync~input .coord_x = 0;
defparam \cam_vsync~input .coord_y = 9;
defparam \cam_vsync~input .coord_z = 2;
defparam \cam_vsync~input .IN_ASYNC_MODE = 1'b0;
defparam \cam_vsync~input .IN_SYNC_MODE = 1'b0;
defparam \cam_vsync~input .IN_POWERUP = 1'b0;
defparam \cam_vsync~input .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_vsync~input .IN_SYNC_DISABLE = 1'b0;
defparam \cam_vsync~input .OUT_REG_MODE = 1'b0;
defparam \cam_vsync~input .OUT_ASYNC_MODE = 1'b0;
defparam \cam_vsync~input .OUT_SYNC_MODE = 1'b0;
defparam \cam_vsync~input .OUT_POWERUP = 1'b0;
defparam \cam_vsync~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_vsync~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_vsync~input .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_vsync~input .OUT_DDIO = 1'b0;
defparam \cam_vsync~input .OE_REG_MODE = 1'b0;
defparam \cam_vsync~input .OE_ASYNC_MODE = 1'b0;
defparam \cam_vsync~input .OE_SYNC_MODE = 1'b0;
defparam \cam_vsync~input .OE_POWERUP = 1'b0;
defparam \cam_vsync~input .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_vsync~input .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_vsync~input .OE_SYNC_DISABLE = 1'b0;
defparam \cam_vsync~input .OE_DDIO = 1'b0;
defparam \cam_vsync~input .CFG_TRI_INPUT = 1'b0;
defparam \cam_vsync~input .CFG_PULL_UP = 1'b0;
defparam \cam_vsync~input .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_vsync~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_vsync~input .CFG_PDRV = 7'b0011010;
defparam \cam_vsync~input .CFG_NDRV = 7'b0011000;
defparam \cam_vsync~input .CFG_KEEP = 2'b00;
defparam \cam_vsync~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_vsync~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_vsync~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_vsync~input .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_vsync~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_vsync~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_vsync~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_vsync~input .CFG_OSCDIV = 2'b00;
defparam \cam_vsync~input .CFG_ROCTUSR = 1'b0;
defparam \cam_vsync~input .CFG_SEL_CUA = 1'b0;
defparam \cam_vsync~input .CFG_ROCT_EN = 1'b0;
defparam \cam_vsync~input .INPUT_ONLY = 1'b0;
defparam \cam_vsync~input .DPCLK_DELAY = 4'b0000;
defparam \cam_vsync~input .OUT_DELAY = 1'b0;
defparam \cam_vsync~input .IN_DATA_DELAY = 3'b000;
defparam \cam_vsync~input .IN_REG_DELAY = 3'b000;

alta_dio \cam_xclk~output (
	.padio(cam_xclk),
	.datain(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \cam_xclk~output .coord_x = 0;
defparam \cam_xclk~output .coord_y = 5;
defparam \cam_xclk~output .coord_z = 0;
defparam \cam_xclk~output .IN_ASYNC_MODE = 1'b0;
defparam \cam_xclk~output .IN_SYNC_MODE = 1'b0;
defparam \cam_xclk~output .IN_POWERUP = 1'b0;
defparam \cam_xclk~output .IN_ASYNC_DISABLE = 1'b0;
defparam \cam_xclk~output .IN_SYNC_DISABLE = 1'b0;
defparam \cam_xclk~output .OUT_REG_MODE = 1'b0;
defparam \cam_xclk~output .OUT_ASYNC_MODE = 1'b0;
defparam \cam_xclk~output .OUT_SYNC_MODE = 1'b0;
defparam \cam_xclk~output .OUT_POWERUP = 1'b0;
defparam \cam_xclk~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \cam_xclk~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \cam_xclk~output .OUT_SYNC_DISABLE = 1'b0;
defparam \cam_xclk~output .OUT_DDIO = 1'b0;
defparam \cam_xclk~output .OE_REG_MODE = 1'b0;
defparam \cam_xclk~output .OE_ASYNC_MODE = 1'b0;
defparam \cam_xclk~output .OE_SYNC_MODE = 1'b0;
defparam \cam_xclk~output .OE_POWERUP = 1'b0;
defparam \cam_xclk~output .OE_CLKEN_DISABLE = 1'b0;
defparam \cam_xclk~output .OE_ASYNC_DISABLE = 1'b0;
defparam \cam_xclk~output .OE_SYNC_DISABLE = 1'b0;
defparam \cam_xclk~output .OE_DDIO = 1'b0;
defparam \cam_xclk~output .CFG_TRI_INPUT = 1'b0;
defparam \cam_xclk~output .CFG_PULL_UP = 1'b0;
defparam \cam_xclk~output .CFG_OPEN_DRAIN = 1'b0;
defparam \cam_xclk~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \cam_xclk~output .CFG_PDRV = 7'b0011010;
defparam \cam_xclk~output .CFG_NDRV = 7'b0011000;
defparam \cam_xclk~output .CFG_KEEP = 2'b00;
defparam \cam_xclk~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \cam_xclk~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \cam_xclk~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \cam_xclk~output .CFG_LVDS_IN_EN = 1'b0;
defparam \cam_xclk~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \cam_xclk~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \cam_xclk~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \cam_xclk~output .CFG_OSCDIV = 2'b00;
defparam \cam_xclk~output .CFG_ROCTUSR = 1'b0;
defparam \cam_xclk~output .CFG_SEL_CUA = 1'b0;
defparam \cam_xclk~output .CFG_ROCT_EN = 1'b0;
defparam \cam_xclk~output .INPUT_ONLY = 1'b0;
defparam \cam_xclk~output .DPCLK_DELAY = 4'b0000;
defparam \cam_xclk~output .OUT_DELAY = 1'b0;
defparam \cam_xclk~output .IN_DATA_DELAY = 3'b000;
defparam \cam_xclk~output .IN_REG_DELAY = 3'b000;

alta_slice \camera_if_inst|Equal0~0 (
	.A(\camera_if_inst|v_cnt [3]),
	.B(\camera_if_inst|v_cnt [2]),
	.C(\camera_if_inst|v_cnt [1]),
	.D(\camera_if_inst|v_cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal0~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal0~0 .coord_x = 6;
defparam \camera_if_inst|Equal0~0 .coord_y = 11;
defparam \camera_if_inst|Equal0~0 .coord_z = 7;
defparam \camera_if_inst|Equal0~0 .mask = 16'hFFFE;
defparam \camera_if_inst|Equal0~0 .modeMux = 1'b0;
defparam \camera_if_inst|Equal0~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal0~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal0~0 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal0~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal0~1 (
	.A(\camera_if_inst|v_cnt [5]),
	.B(\camera_if_inst|v_cnt [6]),
	.C(\camera_if_inst|v_cnt [4]),
	.D(\camera_if_inst|v_cnt [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal0~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal0~1 .coord_x = 11;
defparam \camera_if_inst|Equal0~1 .coord_y = 11;
defparam \camera_if_inst|Equal0~1 .coord_z = 3;
defparam \camera_if_inst|Equal0~1 .mask = 16'hFFFE;
defparam \camera_if_inst|Equal0~1 .modeMux = 1'b0;
defparam \camera_if_inst|Equal0~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal0~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal0~1 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal0~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal0~2 (
	.A(\camera_if_inst|v_cnt [9]),
	.B(\camera_if_inst|v_cnt [8]),
	.C(\camera_if_inst|v_cnt [10]),
	.D(\camera_if_inst|v_cnt [11]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal0~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal0~2 .coord_x = 9;
defparam \camera_if_inst|Equal0~2 .coord_y = 11;
defparam \camera_if_inst|Equal0~2 .coord_z = 7;
defparam \camera_if_inst|Equal0~2 .mask = 16'hFFFE;
defparam \camera_if_inst|Equal0~2 .modeMux = 1'b0;
defparam \camera_if_inst|Equal0~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal0~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal0~2 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal0~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal0~3 (
	.A(\camera_if_inst|v_cnt [15]),
	.B(\camera_if_inst|v_cnt [14]),
	.C(\camera_if_inst|v_cnt [12]),
	.D(\camera_if_inst|v_cnt [13]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal0~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal0~3 .coord_x = 7;
defparam \camera_if_inst|Equal0~3 .coord_y = 11;
defparam \camera_if_inst|Equal0~3 .coord_z = 15;
defparam \camera_if_inst|Equal0~3 .mask = 16'hFFFE;
defparam \camera_if_inst|Equal0~3 .modeMux = 1'b0;
defparam \camera_if_inst|Equal0~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal0~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal0~3 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal0~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal0~4 (
	.A(\camera_if_inst|Equal0~3_combout ),
	.B(\camera_if_inst|Equal0~1_combout ),
	.C(\camera_if_inst|Equal0~2_combout ),
	.D(\camera_if_inst|Equal0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal0~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal0~4 .coord_x = 10;
defparam \camera_if_inst|Equal0~4 .coord_y = 11;
defparam \camera_if_inst|Equal0~4 .coord_z = 10;
defparam \camera_if_inst|Equal0~4 .mask = 16'hFFFE;
defparam \camera_if_inst|Equal0~4 .modeMux = 1'b0;
defparam \camera_if_inst|Equal0~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal0~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal0~4 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal0~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal2~0 (
	.A(\camera_if_inst|f_cnt [1]),
	.B(\camera_if_inst|f_cnt [2]),
	.C(vcc),
	.D(\camera_if_inst|f_cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal2~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal2~0 .coord_x = 5;
defparam \camera_if_inst|Equal2~0 .coord_y = 11;
defparam \camera_if_inst|Equal2~0 .coord_z = 4;
defparam \camera_if_inst|Equal2~0 .mask = 16'h8800;
defparam \camera_if_inst|Equal2~0 .modeMux = 1'b0;
defparam \camera_if_inst|Equal2~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal2~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal2~0 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal2~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal3~0 (
	.A(\camera_if_inst|h_cnt [1]),
	.B(\camera_if_inst|h_cnt [3]),
	.C(\camera_if_inst|h_cnt [2]),
	.D(\camera_if_inst|h_cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal3~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal3~0 .coord_x = 5;
defparam \camera_if_inst|Equal3~0 .coord_y = 11;
defparam \camera_if_inst|Equal3~0 .coord_z = 8;
defparam \camera_if_inst|Equal3~0 .mask = 16'h7FFF;
defparam \camera_if_inst|Equal3~0 .modeMux = 1'b0;
defparam \camera_if_inst|Equal3~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal3~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal3~0 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal3~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal3~1 (
	.A(\camera_if_inst|h_cnt [6]),
	.B(\camera_if_inst|h_cnt [5]),
	.C(\camera_if_inst|h_cnt [7]),
	.D(\camera_if_inst|h_cnt [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal3~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal3~1 .coord_x = 5;
defparam \camera_if_inst|Equal3~1 .coord_y = 11;
defparam \camera_if_inst|Equal3~1 .coord_z = 9;
defparam \camera_if_inst|Equal3~1 .mask = 16'hF7FF;
defparam \camera_if_inst|Equal3~1 .modeMux = 1'b0;
defparam \camera_if_inst|Equal3~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal3~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal3~1 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal3~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal3~2 (
	.A(vcc),
	.B(\camera_if_inst|Equal3~0_combout ),
	.C(vcc),
	.D(\camera_if_inst|Equal3~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal3~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal3~2 .coord_x = 5;
defparam \camera_if_inst|Equal3~2 .coord_y = 11;
defparam \camera_if_inst|Equal3~2 .coord_z = 13;
defparam \camera_if_inst|Equal3~2 .mask = 16'hFFCC;
defparam \camera_if_inst|Equal3~2 .modeMux = 1'b0;
defparam \camera_if_inst|Equal3~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal3~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal3~2 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal3~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal3~3 (
	.A(\camera_if_inst|h_cnt [8]),
	.B(\camera_if_inst|h_cnt [11]),
	.C(\camera_if_inst|h_cnt [9]),
	.D(\camera_if_inst|h_cnt [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal3~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal3~3 .coord_x = 5;
defparam \camera_if_inst|Equal3~3 .coord_y = 11;
defparam \camera_if_inst|Equal3~3 .coord_z = 5;
defparam \camera_if_inst|Equal3~3 .mask = 16'hFFEF;
defparam \camera_if_inst|Equal3~3 .modeMux = 1'b0;
defparam \camera_if_inst|Equal3~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal3~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal3~3 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal3~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|Equal3~4 (
	.A(\camera_if_inst|h_cnt [15]),
	.B(\camera_if_inst|h_cnt [13]),
	.C(\camera_if_inst|h_cnt [14]),
	.D(\camera_if_inst|h_cnt [12]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|Equal3~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|Equal3~4 .coord_x = 5;
defparam \camera_if_inst|Equal3~4 .coord_y = 11;
defparam \camera_if_inst|Equal3~4 .coord_z = 10;
defparam \camera_if_inst|Equal3~4 .mask = 16'hFFFE;
defparam \camera_if_inst|Equal3~4 .modeMux = 1'b0;
defparam \camera_if_inst|Equal3~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|Equal3~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|Equal3~4 .BypassEn = 1'b0;
defparam \camera_if_inst|Equal3~4 .CarryEnb = 1'b1;

alta_io_gclk \camera_if_inst|Equal4~0clkctrl (
	.inclk(\camera_if_inst|Equal4~0_combout ),
	.outclk(\camera_if_inst|Equal4~0clkctrl_outclk ));
defparam \camera_if_inst|Equal4~0clkctrl .coord_x = 0;
defparam \camera_if_inst|Equal4~0clkctrl .coord_y = 12;
defparam \camera_if_inst|Equal4~0clkctrl .coord_z = 4;

alta_slice \camera_if_inst|cam_data_r0[0] (
	.A(),
	.B(),
	.C(\cam_data[0]~input_o ),
	.D(),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [0]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(SyncReset_X9_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X9_Y7_VCC),
	.LutOut(),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [0]));
defparam \camera_if_inst|cam_data_r0[0] .coord_x = 10;
defparam \camera_if_inst|cam_data_r0[0] .coord_y = 11;
defparam \camera_if_inst|cam_data_r0[0] .coord_z = 15;
defparam \camera_if_inst|cam_data_r0[0] .mask = 16'hFFFF;
defparam \camera_if_inst|cam_data_r0[0] .modeMux = 1'b1;
defparam \camera_if_inst|cam_data_r0[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[0] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_data_r0[0] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[1] (
	.A(),
	.B(),
	.C(\cam_data[1]~input_o ),
	.D(),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [1]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(SyncReset_X9_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X9_Y7_VCC),
	.LutOut(),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [1]));
defparam \camera_if_inst|cam_data_r0[1] .coord_x = 10;
defparam \camera_if_inst|cam_data_r0[1] .coord_y = 11;
defparam \camera_if_inst|cam_data_r0[1] .coord_z = 11;
defparam \camera_if_inst|cam_data_r0[1] .mask = 16'hFFFF;
defparam \camera_if_inst|cam_data_r0[1] .modeMux = 1'b1;
defparam \camera_if_inst|cam_data_r0[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[1] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_data_r0[1] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[2] (
	.A(),
	.B(),
	.C(\cam_data[2]~input_o ),
	.D(),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [2]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(SyncReset_X9_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X9_Y7_VCC),
	.LutOut(),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [2]));
defparam \camera_if_inst|cam_data_r0[2] .coord_x = 10;
defparam \camera_if_inst|cam_data_r0[2] .coord_y = 11;
defparam \camera_if_inst|cam_data_r0[2] .coord_z = 7;
defparam \camera_if_inst|cam_data_r0[2] .mask = 16'hFFFF;
defparam \camera_if_inst|cam_data_r0[2] .modeMux = 1'b1;
defparam \camera_if_inst|cam_data_r0[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[2] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_data_r0[2] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[3] (
	.A(\camera_if_inst|cam_data_r0 [1]),
	.B(\camera_if_inst|cam_data_r0 [2]),
	.C(\cam_data[3]~input_o ),
	.D(\camera_if_inst|cam_data_r0 [0]),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [3]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(SyncReset_X9_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X9_Y7_VCC),
	.LutOut(\camera_if_inst|Equal1~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [3]));
defparam \camera_if_inst|cam_data_r0[3] .coord_x = 10;
defparam \camera_if_inst|cam_data_r0[3] .coord_y = 11;
defparam \camera_if_inst|cam_data_r0[3] .coord_z = 0;
defparam \camera_if_inst|cam_data_r0[3] .mask = 16'hFFFE;
defparam \camera_if_inst|cam_data_r0[3] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[3] .FeedbackMux = 1'b1;
defparam \camera_if_inst|cam_data_r0[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[3] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_data_r0[3] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cam_data[4]~input_o ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [4]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r0[4]~feeder_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [4]));
defparam \camera_if_inst|cam_data_r0[4] .coord_x = 10;
defparam \camera_if_inst|cam_data_r0[4] .coord_y = 11;
defparam \camera_if_inst|cam_data_r0[4] .coord_z = 3;
defparam \camera_if_inst|cam_data_r0[4] .mask = 16'hFF00;
defparam \camera_if_inst|cam_data_r0[4] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[4] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r0[4] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[5] (
	.A(\camera_if_inst|cam_data_r0 [4]),
	.B(\camera_if_inst|cam_data_r0 [6]),
	.C(\cam_data[5]~input_o ),
	.D(\camera_if_inst|cam_data_r0 [7]),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [5]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(SyncReset_X9_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X9_Y7_VCC),
	.LutOut(\camera_if_inst|Equal1~1_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [5]));
defparam \camera_if_inst|cam_data_r0[5] .coord_x = 10;
defparam \camera_if_inst|cam_data_r0[5] .coord_y = 11;
defparam \camera_if_inst|cam_data_r0[5] .coord_z = 14;
defparam \camera_if_inst|cam_data_r0[5] .mask = 16'hFFFE;
defparam \camera_if_inst|cam_data_r0[5] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[5] .FeedbackMux = 1'b1;
defparam \camera_if_inst|cam_data_r0[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[5] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_data_r0[5] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[6] (
	.A(),
	.B(),
	.C(\cam_data[6]~input_o ),
	.D(),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [6]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(SyncReset_X9_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X9_Y7_VCC),
	.LutOut(),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [6]));
defparam \camera_if_inst|cam_data_r0[6] .coord_x = 10;
defparam \camera_if_inst|cam_data_r0[6] .coord_y = 11;
defparam \camera_if_inst|cam_data_r0[6] .coord_z = 12;
defparam \camera_if_inst|cam_data_r0[6] .mask = 16'hFFFF;
defparam \camera_if_inst|cam_data_r0[6] .modeMux = 1'b1;
defparam \camera_if_inst|cam_data_r0[6] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[6] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[6] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_data_r0[6] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r0[7] (
	.A(),
	.B(),
	.C(\cam_data[7]~input_o ),
	.D(),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r0 [7]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(SyncReset_X2_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_VCC),
	.LutOut(),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r0 [7]));
defparam \camera_if_inst|cam_data_r0[7] .coord_x = 5;
defparam \camera_if_inst|cam_data_r0[7] .coord_y = 11;
defparam \camera_if_inst|cam_data_r0[7] .coord_z = 0;
defparam \camera_if_inst|cam_data_r0[7] .mask = 16'hFFFF;
defparam \camera_if_inst|cam_data_r0[7] .modeMux = 1'b1;
defparam \camera_if_inst|cam_data_r0[7] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[7] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r0[7] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_data_r0[7] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[0] (
	.A(\camera_if_inst|Equal0~4_combout ),
	.B(\camera_if_inst|cam_data_r0 [0]),
	.C(\camera_if_inst|Equal1~0_combout ),
	.D(\camera_if_inst|Equal1~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [0]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~6_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [0]));
defparam \camera_if_inst|cam_data_r1[0] .coord_x = 10;
defparam \camera_if_inst|cam_data_r1[0] .coord_y = 11;
defparam \camera_if_inst|cam_data_r1[0] .coord_z = 8;
defparam \camera_if_inst|cam_data_r1[0] .mask = 16'h888A;
defparam \camera_if_inst|cam_data_r1[0] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[0] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[0] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[1] (
	.A(\camera_if_inst|cam_data_r0 [1]),
	.B(\camera_if_inst|Equal0~4_combout ),
	.C(\camera_if_inst|Equal1~0_combout ),
	.D(\camera_if_inst|Equal1~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [1]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~4_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [1]));
defparam \camera_if_inst|cam_data_r1[1] .coord_x = 10;
defparam \camera_if_inst|cam_data_r1[1] .coord_y = 11;
defparam \camera_if_inst|cam_data_r1[1] .coord_z = 9;
defparam \camera_if_inst|cam_data_r1[1] .mask = 16'h8880;
defparam \camera_if_inst|cam_data_r1[1] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[1] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[1] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[2] (
	.A(\camera_if_inst|Equal0~4_combout ),
	.B(\camera_if_inst|cam_data_r0 [2]),
	.C(\camera_if_inst|Equal1~0_combout ),
	.D(\camera_if_inst|Equal1~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [2]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~3_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [2]));
defparam \camera_if_inst|cam_data_r1[2] .coord_x = 10;
defparam \camera_if_inst|cam_data_r1[2] .coord_y = 11;
defparam \camera_if_inst|cam_data_r1[2] .coord_z = 13;
defparam \camera_if_inst|cam_data_r1[2] .mask = 16'h8880;
defparam \camera_if_inst|cam_data_r1[2] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[2] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[2] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[3] (
	.A(\camera_if_inst|cam_data_r0 [3]),
	.B(\camera_if_inst|Equal0~4_combout ),
	.C(\camera_if_inst|Equal1~0_combout ),
	.D(\camera_if_inst|Equal1~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [3]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~5_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [3]));
defparam \camera_if_inst|cam_data_r1[3] .coord_x = 10;
defparam \camera_if_inst|cam_data_r1[3] .coord_y = 11;
defparam \camera_if_inst|cam_data_r1[3] .coord_z = 5;
defparam \camera_if_inst|cam_data_r1[3] .mask = 16'h8880;
defparam \camera_if_inst|cam_data_r1[3] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[3] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[3] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[3] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[4] (
	.A(\camera_if_inst|cam_data_r0 [4]),
	.B(\camera_if_inst|Equal0~4_combout ),
	.C(\camera_if_inst|Equal1~0_combout ),
	.D(\camera_if_inst|Equal1~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [4]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~7_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [4]));
defparam \camera_if_inst|cam_data_r1[4] .coord_x = 10;
defparam \camera_if_inst|cam_data_r1[4] .coord_y = 11;
defparam \camera_if_inst|cam_data_r1[4] .coord_z = 2;
defparam \camera_if_inst|cam_data_r1[4] .mask = 16'h8880;
defparam \camera_if_inst|cam_data_r1[4] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[4] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[4] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[5] (
	.A(\camera_if_inst|cam_data_r0 [5]),
	.B(\camera_if_inst|Equal0~4_combout ),
	.C(\camera_if_inst|Equal1~0_combout ),
	.D(\camera_if_inst|Equal1~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [5]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [5]));
defparam \camera_if_inst|cam_data_r1[5] .coord_x = 10;
defparam \camera_if_inst|cam_data_r1[5] .coord_y = 11;
defparam \camera_if_inst|cam_data_r1[5] .coord_z = 6;
defparam \camera_if_inst|cam_data_r1[5] .mask = 16'h8880;
defparam \camera_if_inst|cam_data_r1[5] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[5] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[5] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[5] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[6] (
	.A(\camera_if_inst|Equal0~4_combout ),
	.B(\camera_if_inst|cam_data_r0 [6]),
	.C(\camera_if_inst|Equal1~0_combout ),
	.D(\camera_if_inst|Equal1~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [6]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [6]));
defparam \camera_if_inst|cam_data_r1[6] .coord_x = 10;
defparam \camera_if_inst|cam_data_r1[6] .coord_y = 11;
defparam \camera_if_inst|cam_data_r1[6] .coord_z = 4;
defparam \camera_if_inst|cam_data_r1[6] .mask = 16'h8880;
defparam \camera_if_inst|cam_data_r1[6] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[6] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[6] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[6] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[6] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_data_r1[7] (
	.A(\camera_if_inst|Equal0~4_combout ),
	.B(\camera_if_inst|cam_data_r0 [7]),
	.C(\camera_if_inst|Equal1~0_combout ),
	.D(\camera_if_inst|Equal1~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|cam_data_r1 [7]),
	.Clk(\cam_pclk~input_o_X9_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X9_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_data_r1~1_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_data_r1 [7]));
defparam \camera_if_inst|cam_data_r1[7] .coord_x = 10;
defparam \camera_if_inst|cam_data_r1[7] .coord_y = 11;
defparam \camera_if_inst|cam_data_r1[7] .coord_z = 1;
defparam \camera_if_inst|cam_data_r1[7] .mask = 16'h8880;
defparam \camera_if_inst|cam_data_r1[7] .modeMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[7] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[7] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_data_r1[7] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_data_r1[7] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_hsync_r[0] (
	.A(\camera_if_inst|f_cnt [3]),
	.B(vcc),
	.C(\camera_if_inst|Equal2~0_combout ),
	.D(\cam_hsync~input_o ),
	.Cin(),
	.Qin(\camera_if_inst|cam_hsync_r [0]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_hsync_r~1_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_hsync_r [0]));
defparam \camera_if_inst|cam_hsync_r[0] .coord_x = 5;
defparam \camera_if_inst|cam_hsync_r[0] .coord_y = 11;
defparam \camera_if_inst|cam_hsync_r[0] .coord_z = 2;
defparam \camera_if_inst|cam_hsync_r[0] .mask = 16'hA000;
defparam \camera_if_inst|cam_hsync_r[0] .modeMux = 1'b0;
defparam \camera_if_inst|cam_hsync_r[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_hsync_r[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_hsync_r[0] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_hsync_r[0] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_hsync_r[1] (
	.A(\camera_if_inst|f_cnt [3]),
	.B(\camera_if_inst|cam_hsync_r [0]),
	.C(\camera_if_inst|Equal2~0_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|cam_hsync_r [1]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|cam_hsync_r~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_hsync_r [1]));
defparam \camera_if_inst|cam_hsync_r[1] .coord_x = 5;
defparam \camera_if_inst|cam_hsync_r[1] .coord_y = 11;
defparam \camera_if_inst|cam_hsync_r[1] .coord_z = 1;
defparam \camera_if_inst|cam_hsync_r[1] .mask = 16'h8080;
defparam \camera_if_inst|cam_hsync_r[1] .modeMux = 1'b0;
defparam \camera_if_inst|cam_hsync_r[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|cam_hsync_r[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_hsync_r[1] .BypassEn = 1'b0;
defparam \camera_if_inst|cam_hsync_r[1] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_vsync_r[0] (
	.A(\camera_if_inst|f_cnt [3]),
	.B(\camera_if_inst|Equal2~0_combout ),
	.C(\cam_vsync~input_o ),
	.D(\camera_if_inst|cam_vsync_r [1]),
	.Cin(),
	.Qin(\camera_if_inst|cam_vsync_r [0]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(SyncReset_X2_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_VCC),
	.LutOut(\camera_if_inst|f_cnt[3]~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_vsync_r [0]));
defparam \camera_if_inst|cam_vsync_r[0] .coord_x = 5;
defparam \camera_if_inst|cam_vsync_r[0] .coord_y = 11;
defparam \camera_if_inst|cam_vsync_r[0] .coord_z = 7;
defparam \camera_if_inst|cam_vsync_r[0] .mask = 16'h0700;
defparam \camera_if_inst|cam_vsync_r[0] .modeMux = 1'b0;
defparam \camera_if_inst|cam_vsync_r[0] .FeedbackMux = 1'b1;
defparam \camera_if_inst|cam_vsync_r[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_vsync_r[0] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_vsync_r[0] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|cam_vsync_r[1] (
	.A(vcc),
	.B(vcc),
	.C(\camera_if_inst|cam_vsync_r [0]),
	.D(\camera_if_inst|cam_vsync_r [0]),
	.Cin(),
	.Qin(\camera_if_inst|cam_vsync_r [1]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(SyncReset_X2_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X2_Y7_VCC),
	.LutOut(\camera_if_inst|Equal4~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|cam_vsync_r [1]));
defparam \camera_if_inst|cam_vsync_r[1] .coord_x = 5;
defparam \camera_if_inst|cam_vsync_r[1] .coord_y = 11;
defparam \camera_if_inst|cam_vsync_r[1] .coord_z = 11;
defparam \camera_if_inst|cam_vsync_r[1] .mask = 16'h00F0;
defparam \camera_if_inst|cam_vsync_r[1] .modeMux = 1'b0;
defparam \camera_if_inst|cam_vsync_r[1] .FeedbackMux = 1'b1;
defparam \camera_if_inst|cam_vsync_r[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|cam_vsync_r[1] .BypassEn = 1'b1;
defparam \camera_if_inst|cam_vsync_r[1] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|f_cnt[0] (
	.A(\camera_if_inst|f_cnt [3]),
	.B(\camera_if_inst|Equal2~0_combout ),
	.C(vcc),
	.D(\camera_if_inst|Equal4~0_combout ),
	.Cin(),
	.Qin(\camera_if_inst|f_cnt [0]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|f_cnt[0]~5_combout ),
	.Cout(),
	.Q(\camera_if_inst|f_cnt [0]));
defparam \camera_if_inst|f_cnt[0] .coord_x = 5;
defparam \camera_if_inst|f_cnt[0] .coord_y = 11;
defparam \camera_if_inst|f_cnt[0] .coord_z = 6;
defparam \camera_if_inst|f_cnt[0] .mask = 16'h87F0;
defparam \camera_if_inst|f_cnt[0] .modeMux = 1'b0;
defparam \camera_if_inst|f_cnt[0] .FeedbackMux = 1'b1;
defparam \camera_if_inst|f_cnt[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|f_cnt[0] .BypassEn = 1'b0;
defparam \camera_if_inst|f_cnt[0] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|f_cnt[1] (
	.A(vcc),
	.B(\camera_if_inst|f_cnt[3]~2_combout ),
	.C(vcc),
	.D(\camera_if_inst|f_cnt [0]),
	.Cin(),
	.Qin(\camera_if_inst|f_cnt [1]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|f_cnt[1]~4_combout ),
	.Cout(),
	.Q(\camera_if_inst|f_cnt [1]));
defparam \camera_if_inst|f_cnt[1] .coord_x = 5;
defparam \camera_if_inst|f_cnt[1] .coord_y = 11;
defparam \camera_if_inst|f_cnt[1] .coord_z = 3;
defparam \camera_if_inst|f_cnt[1] .mask = 16'h3CF0;
defparam \camera_if_inst|f_cnt[1] .modeMux = 1'b0;
defparam \camera_if_inst|f_cnt[1] .FeedbackMux = 1'b1;
defparam \camera_if_inst|f_cnt[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|f_cnt[1] .BypassEn = 1'b0;
defparam \camera_if_inst|f_cnt[1] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|f_cnt[2] (
	.A(\camera_if_inst|f_cnt [1]),
	.B(\camera_if_inst|f_cnt[3]~2_combout ),
	.C(vcc),
	.D(\camera_if_inst|f_cnt [0]),
	.Cin(),
	.Qin(\camera_if_inst|f_cnt [2]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|f_cnt[2]~3_combout ),
	.Cout(),
	.Q(\camera_if_inst|f_cnt [2]));
defparam \camera_if_inst|f_cnt[2] .coord_x = 5;
defparam \camera_if_inst|f_cnt[2] .coord_y = 11;
defparam \camera_if_inst|f_cnt[2] .coord_z = 12;
defparam \camera_if_inst|f_cnt[2] .mask = 16'h78F0;
defparam \camera_if_inst|f_cnt[2] .modeMux = 1'b0;
defparam \camera_if_inst|f_cnt[2] .FeedbackMux = 1'b1;
defparam \camera_if_inst|f_cnt[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|f_cnt[2] .BypassEn = 1'b0;
defparam \camera_if_inst|f_cnt[2] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|f_cnt[3] (
	.A(\camera_if_inst|cam_vsync_r [1]),
	.B(\camera_if_inst|Equal2~0_combout ),
	.C(vcc),
	.D(\camera_if_inst|cam_vsync_r [0]),
	.Cin(),
	.Qin(\camera_if_inst|f_cnt [3]),
	.Clk(\cam_pclk~input_o_X2_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X2_Y7_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|f_cnt[3]~6_combout ),
	.Cout(),
	.Q(\camera_if_inst|f_cnt [3]));
defparam \camera_if_inst|f_cnt[3] .coord_x = 5;
defparam \camera_if_inst|f_cnt[3] .coord_y = 11;
defparam \camera_if_inst|f_cnt[3] .coord_z = 15;
defparam \camera_if_inst|f_cnt[3] .mask = 16'hF0F8;
defparam \camera_if_inst|f_cnt[3] .modeMux = 1'b0;
defparam \camera_if_inst|f_cnt[3] .FeedbackMux = 1'b1;
defparam \camera_if_inst|f_cnt[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|f_cnt[3] .BypassEn = 1'b0;
defparam \camera_if_inst|f_cnt[3] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|h_cnt[0] (
	.A(\camera_if_inst|h_cnt [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|h_cnt [0]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[0]~16_combout ),
	.Cout(\camera_if_inst|h_cnt[0]~17 ),
	.Q(\camera_if_inst|h_cnt [0]));
defparam \camera_if_inst|h_cnt[0] .coord_x = 4;
defparam \camera_if_inst|h_cnt[0] .coord_y = 11;
defparam \camera_if_inst|h_cnt[0] .coord_z = 0;
defparam \camera_if_inst|h_cnt[0] .mask = 16'h55AA;
defparam \camera_if_inst|h_cnt[0] .modeMux = 1'b0;
defparam \camera_if_inst|h_cnt[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[0] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[0] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[10] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [10]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[9]~35 ),
	.Qin(\camera_if_inst|h_cnt [10]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[10]~36_combout ),
	.Cout(\camera_if_inst|h_cnt[10]~37 ),
	.Q(\camera_if_inst|h_cnt [10]));
defparam \camera_if_inst|h_cnt[10] .coord_x = 4;
defparam \camera_if_inst|h_cnt[10] .coord_y = 11;
defparam \camera_if_inst|h_cnt[10] .coord_z = 10;
defparam \camera_if_inst|h_cnt[10] .mask = 16'hC30C;
defparam \camera_if_inst|h_cnt[10] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[10] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[10] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[10] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[10] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[11] (
	.A(\camera_if_inst|h_cnt [11]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[10]~37 ),
	.Qin(\camera_if_inst|h_cnt [11]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[11]~38_combout ),
	.Cout(\camera_if_inst|h_cnt[11]~39 ),
	.Q(\camera_if_inst|h_cnt [11]));
defparam \camera_if_inst|h_cnt[11] .coord_x = 4;
defparam \camera_if_inst|h_cnt[11] .coord_y = 11;
defparam \camera_if_inst|h_cnt[11] .coord_z = 11;
defparam \camera_if_inst|h_cnt[11] .mask = 16'h5A5F;
defparam \camera_if_inst|h_cnt[11] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[11] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[11] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[11] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[11] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[12] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [12]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[11]~39 ),
	.Qin(\camera_if_inst|h_cnt [12]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[12]~40_combout ),
	.Cout(\camera_if_inst|h_cnt[12]~41 ),
	.Q(\camera_if_inst|h_cnt [12]));
defparam \camera_if_inst|h_cnt[12] .coord_x = 4;
defparam \camera_if_inst|h_cnt[12] .coord_y = 11;
defparam \camera_if_inst|h_cnt[12] .coord_z = 12;
defparam \camera_if_inst|h_cnt[12] .mask = 16'hC30C;
defparam \camera_if_inst|h_cnt[12] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[12] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[12] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[12] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[12] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[13] (
	.A(\camera_if_inst|h_cnt [13]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[12]~41 ),
	.Qin(\camera_if_inst|h_cnt [13]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[13]~42_combout ),
	.Cout(\camera_if_inst|h_cnt[13]~43 ),
	.Q(\camera_if_inst|h_cnt [13]));
defparam \camera_if_inst|h_cnt[13] .coord_x = 4;
defparam \camera_if_inst|h_cnt[13] .coord_y = 11;
defparam \camera_if_inst|h_cnt[13] .coord_z = 13;
defparam \camera_if_inst|h_cnt[13] .mask = 16'h5A5F;
defparam \camera_if_inst|h_cnt[13] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[13] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[13] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[13] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[13] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[14] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [14]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[13]~43 ),
	.Qin(\camera_if_inst|h_cnt [14]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[14]~44_combout ),
	.Cout(\camera_if_inst|h_cnt[14]~45 ),
	.Q(\camera_if_inst|h_cnt [14]));
defparam \camera_if_inst|h_cnt[14] .coord_x = 4;
defparam \camera_if_inst|h_cnt[14] .coord_y = 11;
defparam \camera_if_inst|h_cnt[14] .coord_z = 14;
defparam \camera_if_inst|h_cnt[14] .mask = 16'hC30C;
defparam \camera_if_inst|h_cnt[14] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[14] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[14] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[14] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[14] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[15] (
	.A(\camera_if_inst|h_cnt [15]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[14]~45 ),
	.Qin(\camera_if_inst|h_cnt [15]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[15]~46_combout ),
	.Cout(),
	.Q(\camera_if_inst|h_cnt [15]));
defparam \camera_if_inst|h_cnt[15] .coord_x = 4;
defparam \camera_if_inst|h_cnt[15] .coord_y = 11;
defparam \camera_if_inst|h_cnt[15] .coord_z = 15;
defparam \camera_if_inst|h_cnt[15] .mask = 16'h5A5A;
defparam \camera_if_inst|h_cnt[15] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[15] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[15] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[15] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[15] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|h_cnt[1] (
	.A(\camera_if_inst|h_cnt [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[0]~17 ),
	.Qin(\camera_if_inst|h_cnt [1]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[1]~18_combout ),
	.Cout(\camera_if_inst|h_cnt[1]~19 ),
	.Q(\camera_if_inst|h_cnt [1]));
defparam \camera_if_inst|h_cnt[1] .coord_x = 4;
defparam \camera_if_inst|h_cnt[1] .coord_y = 11;
defparam \camera_if_inst|h_cnt[1] .coord_z = 1;
defparam \camera_if_inst|h_cnt[1] .mask = 16'h5A5F;
defparam \camera_if_inst|h_cnt[1] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[1] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[1] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[2] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[1]~19 ),
	.Qin(\camera_if_inst|h_cnt [2]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[2]~20_combout ),
	.Cout(\camera_if_inst|h_cnt[2]~21 ),
	.Q(\camera_if_inst|h_cnt [2]));
defparam \camera_if_inst|h_cnt[2] .coord_x = 4;
defparam \camera_if_inst|h_cnt[2] .coord_y = 11;
defparam \camera_if_inst|h_cnt[2] .coord_z = 2;
defparam \camera_if_inst|h_cnt[2] .mask = 16'hC30C;
defparam \camera_if_inst|h_cnt[2] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[2] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[2] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[3] (
	.A(\camera_if_inst|h_cnt [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[2]~21 ),
	.Qin(\camera_if_inst|h_cnt [3]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[3]~22_combout ),
	.Cout(\camera_if_inst|h_cnt[3]~23 ),
	.Q(\camera_if_inst|h_cnt [3]));
defparam \camera_if_inst|h_cnt[3] .coord_x = 4;
defparam \camera_if_inst|h_cnt[3] .coord_y = 11;
defparam \camera_if_inst|h_cnt[3] .coord_z = 3;
defparam \camera_if_inst|h_cnt[3] .mask = 16'h5A5F;
defparam \camera_if_inst|h_cnt[3] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[3] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[3] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[3] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[4] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[3]~23 ),
	.Qin(\camera_if_inst|h_cnt [4]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[4]~24_combout ),
	.Cout(\camera_if_inst|h_cnt[4]~25 ),
	.Q(\camera_if_inst|h_cnt [4]));
defparam \camera_if_inst|h_cnt[4] .coord_x = 4;
defparam \camera_if_inst|h_cnt[4] .coord_y = 11;
defparam \camera_if_inst|h_cnt[4] .coord_z = 4;
defparam \camera_if_inst|h_cnt[4] .mask = 16'hC30C;
defparam \camera_if_inst|h_cnt[4] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[4] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[4] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[5] (
	.A(\camera_if_inst|h_cnt [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[4]~25 ),
	.Qin(\camera_if_inst|h_cnt [5]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[5]~26_combout ),
	.Cout(\camera_if_inst|h_cnt[5]~27 ),
	.Q(\camera_if_inst|h_cnt [5]));
defparam \camera_if_inst|h_cnt[5] .coord_x = 4;
defparam \camera_if_inst|h_cnt[5] .coord_y = 11;
defparam \camera_if_inst|h_cnt[5] .coord_z = 5;
defparam \camera_if_inst|h_cnt[5] .mask = 16'h5A5F;
defparam \camera_if_inst|h_cnt[5] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[5] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[5] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[5] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[6] (
	.A(\camera_if_inst|h_cnt [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[5]~27 ),
	.Qin(\camera_if_inst|h_cnt [6]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[6]~28_combout ),
	.Cout(\camera_if_inst|h_cnt[6]~29 ),
	.Q(\camera_if_inst|h_cnt [6]));
defparam \camera_if_inst|h_cnt[6] .coord_x = 4;
defparam \camera_if_inst|h_cnt[6] .coord_y = 11;
defparam \camera_if_inst|h_cnt[6] .coord_z = 6;
defparam \camera_if_inst|h_cnt[6] .mask = 16'hA50A;
defparam \camera_if_inst|h_cnt[6] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[6] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[6] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[6] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[6] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[7] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[6]~29 ),
	.Qin(\camera_if_inst|h_cnt [7]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[7]~30_combout ),
	.Cout(\camera_if_inst|h_cnt[7]~31 ),
	.Q(\camera_if_inst|h_cnt [7]));
defparam \camera_if_inst|h_cnt[7] .coord_x = 4;
defparam \camera_if_inst|h_cnt[7] .coord_y = 11;
defparam \camera_if_inst|h_cnt[7] .coord_z = 7;
defparam \camera_if_inst|h_cnt[7] .mask = 16'h3C3F;
defparam \camera_if_inst|h_cnt[7] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[7] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[7] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[7] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[7] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[8] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [8]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[7]~31 ),
	.Qin(\camera_if_inst|h_cnt [8]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[8]~32_combout ),
	.Cout(\camera_if_inst|h_cnt[8]~33 ),
	.Q(\camera_if_inst|h_cnt [8]));
defparam \camera_if_inst|h_cnt[8] .coord_x = 4;
defparam \camera_if_inst|h_cnt[8] .coord_y = 11;
defparam \camera_if_inst|h_cnt[8] .coord_z = 8;
defparam \camera_if_inst|h_cnt[8] .mask = 16'hC30C;
defparam \camera_if_inst|h_cnt[8] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[8] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[8] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[8] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[8] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|h_cnt[9] (
	.A(vcc),
	.B(\camera_if_inst|h_cnt [9]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|h_cnt[8]~33 ),
	.Qin(\camera_if_inst|h_cnt [9]),
	.Clk(\cam_pclk~input_o_X1_Y7_SIG_VCC ),
	.AsyncReset(AsyncReset_X1_Y7_GND),
	.SyncReset(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X1_Y7_GND),
	.LutOut(\camera_if_inst|h_cnt[9]~34_combout ),
	.Cout(\camera_if_inst|h_cnt[9]~35 ),
	.Q(\camera_if_inst|h_cnt [9]));
defparam \camera_if_inst|h_cnt[9] .coord_x = 4;
defparam \camera_if_inst|h_cnt[9] .coord_y = 11;
defparam \camera_if_inst|h_cnt[9] .coord_z = 9;
defparam \camera_if_inst|h_cnt[9] .mask = 16'h3C3F;
defparam \camera_if_inst|h_cnt[9] .modeMux = 1'b1;
defparam \camera_if_inst|h_cnt[9] .FeedbackMux = 1'b0;
defparam \camera_if_inst|h_cnt[9] .ShiftMux = 1'b0;
defparam \camera_if_inst|h_cnt[9] .BypassEn = 1'b1;
defparam \camera_if_inst|h_cnt[9] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] (
	.A(\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.10~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X17_Y11_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0]~22_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .mask = 16'h78F0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .FeedbackMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[0] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1]~7_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1]~8 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .mask = 16'h6688;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[1]~8 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2]~9_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2]~10 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .mask = 16'h3C3F;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[2]~10 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3]~11_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3]~12 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[3]~12 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4]~14_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4]~15 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .mask = 16'h3C3F;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[4]~15 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5]~16_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5]~17 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .mask = 16'hA50A;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[5]~17 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6]~18_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6]~19 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .mask = 16'h3C3F;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[6]~19 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~20_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]));
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .mask = 16'hA5A5;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.B(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.10~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|LessThan1~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .mask = 16'hC400;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan0~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [11]),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [14]),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [13]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [12]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan0~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .mask = 16'h0001;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan0~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan0~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .mask = 16'h0001;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan0~2 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan0~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .mask = 16'h3FFF;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan0~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LessThan0~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [8]),
	.C(\camera_if_inst|u_I2C_AV_Config|LessThan0~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [9]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan0~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .mask = 16'h0032;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan0~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [15]),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [10]),
	.C(\camera_if_inst|u_I2C_AV_Config|LessThan0~3_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LessThan0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .mask = 16'h5100;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan0~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan1~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan1~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .mask = 16'h010F;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|LessThan1~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|LessThan1~0_combout ),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .mask = 16'hF5F5;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|LessThan1~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|Selector3~0 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|Selector3~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .mask = 16'h0C00;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|Selector3~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|Selector3~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .mask = 16'hFFFE;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|Selector3~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|Selector3~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|Selector3~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .mask = 16'hFFFE;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|Selector3~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X28_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~feeder_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~q ));
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .mask = 16'hAAAA;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 (
	.A(\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~q ),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|i2c_en_r0~q ),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|i2c_en_r1~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X28_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y9_SIG ),
	.SyncReset(SyncReset_X28_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X28_Y9_VCC),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|i2c_en_r1~q ));
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .mask = 16'h5050;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .FeedbackMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|i2c_en_r1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [0]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0]~16_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0]~17 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [0]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .mask = 16'h55AA;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [10]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9]~35 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [10]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10]~36_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10]~37 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [10]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [11]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[10]~37 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [11]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11]~38_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11]~39 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [11]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [12]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[11]~39 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [12]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12]~40_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12]~41 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [12]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [13]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[12]~41 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [13]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13]~42_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13]~43 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [13]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [14]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[13]~43 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [14]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14]~44_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14]~45 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [14]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [15]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[14]~45 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [15]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15]~46_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [15]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .mask = 16'h5A5A;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[15] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[0]~17 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [1]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1]~18_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1]~19 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [1]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[1]~19 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [2]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2]~20_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2]~21 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [2]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[2]~21 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [3]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3]~22_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3]~23 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [3]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[3]~23 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [4]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4]~24_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4]~25 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [4]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[4]~25 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [5]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5]~26_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5]~27 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [5]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .mask = 16'h5A5F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[5]~27 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [6]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6]~28_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6]~29 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [6]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .mask = 16'hA50A;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[6]~29 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [7]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7]~30_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7]~31 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [7]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .mask = 16'h3C3F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [8]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[7]~31 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [8]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8]~32_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8]~33 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [8]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [9]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[8]~33 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [9]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X29_Y9_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X29_Y9_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9]~34_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9]~35 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV [9]));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .mask = 16'h3C3F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CLK_DIV[9] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X28_Y9_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X28_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~q ));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .mask = 16'hF00F;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .FeedbackMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_GO (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.00~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~1_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .mask = 16'hB030;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.B(vcc),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .mask = 16'h5500;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_GO~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mI2C_WR (
	.A(\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|Selector3~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.00~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|Selector3~2_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ));
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .mask = 16'h8A88;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mI2C_WR .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 (
	.A(\camera_if_inst|u_I2C_AV_Config|mSetup_ST~11_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACK~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.00~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mSetup_ST~12_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.00~q ));
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .mask = 16'h1500;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.00 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|LessThan1~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.10~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mSetup_ST~10_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ));
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .mask = 16'h0031;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.01 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACK~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|LessThan1~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.10~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X16_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mSetup_ST~13_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.10~q ));
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .mask = 16'h4000;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST.10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 (
	.A(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.00~q ),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|mSetup_ST.01~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|mSetup_ST~11_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .mask = 16'h0F0A;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|mSetup_ST~11 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .mask = 16'h40C0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\cam_sda~input_o ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .mask = 16'h08A8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Selector9~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .mask = 16'hCCD8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR1~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .mask = 16'h0070;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(\cam_sda~input_o ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .mask = 16'h005D;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|END~2_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Selector8~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .mask = 16'h0AFB;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR2~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~3_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .mask = 16'h002A;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 (
	.A(vcc),
	.B(\cam_sda~input_o ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .mask = 16'hCF0F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .mask = 16'h8008;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .mask = 16'hF313;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKR3~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .mask = 16'h3010;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\cam_sda~input_o ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .mask = 16'hD500;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Selector9~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|END~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .mask = 16'h7475;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW1~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .mask = 16'hC040;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~q ),
	.B(\cam_sda~input_o ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .mask = 16'hA030;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Selector8~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .mask = 16'hACAA;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW2~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y11_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~2_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .mask = 16'h2300;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(\cam_sda~input_o ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .mask = 16'hC444;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Selector2~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|END~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .mask = 16'h7475;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACKW3~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKR2~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKR1~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACKR3~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACK~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .mask = 16'h007F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|ACKW1~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|ACKW2~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACKW3~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACK~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .mask = 16'h7F00;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 (
	.A(vcc),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|ACK~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|ACK~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|ACK~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .mask = 16'hFFF0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|ACK~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .mask = 16'h0033;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 (
	.A(vcc),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .mask = 16'h000F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .mask = 16'h0400;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Decoder0~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|END~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|END~5_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y10_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~6_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|END~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .mask = 16'hE0A0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(vcc),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .mask = 16'hAA00;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|END~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .mask = 16'hAA2A;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END~2 (
	.A(vcc),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .mask = 16'h000F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|END~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .mask = 16'h8000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END~4 (
	.A(vcc),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .mask = 16'hF000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|END~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|END~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|END~3_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|END~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|END~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .mask = 16'hF8F0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|END~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .mask = 16'h0033;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .mask = 16'h8000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal0~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Equal3~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .mask = 16'h0004;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Equal3~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Equal3~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .mask = 16'hC000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal3~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Equal5~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .mask = 16'h0080;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Equal5~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~29_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~10_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y10_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X17_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~0_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .mask = 16'h04C4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .mask = 16'hEAC0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|comb~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .mask = 16'h7520;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_CTRL_CLK~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .mask = 16'hD155;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Equal3~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .mask = 16'hCCFA;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .mask = 16'h00DC;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .mask = 16'h1000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~3_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .mask = 16'h0504;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .mask = 16'h2664;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .mask = 16'hCCA8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~7_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .mask = 16'hF3BC;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~5_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~8_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .mask = 16'hFFAE;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|I2C_SCLK~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 (
	.A(vcc),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .mask = 16'hF000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .mask = 16'h0033;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~9_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~7_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .mask = 16'hFFF8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~11_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .mask = 16'h3055;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~11 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~11_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~12_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .mask = 16'h9810;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~12 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~13_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .mask = 16'hFA44;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~13 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~13_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~14_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .mask = 16'hF588;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~14 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|comb~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~15_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .mask = 16'hD800;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~15 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~16_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .mask = 16'h88A0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~16 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~17_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .mask = 16'h5044;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~17 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~15_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~17_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~16_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~18_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .mask = 16'hBBBA;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~18 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~18_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~14_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~19_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .mask = 16'h7520;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~19 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .mask = 16'h0102;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~20_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .mask = 16'h3703;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~20 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~20_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~19_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~21_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .mask = 16'hAEA4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~21 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~22_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .mask = 16'h4450;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~22 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~23_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .mask = 16'hA808;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~23 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~24_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .mask = 16'h0AFA;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~24 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~24_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~25_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .mask = 16'hAEA3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~25 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~26_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .mask = 16'hBA98;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~26 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~26_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~27_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .mask = 16'hF588;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~27 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~27_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~31_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~25_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~28_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .mask = 16'hDDA0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~28 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~28_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~12_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~21_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~29_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .mask = 16'hDDA0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~29 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .mask = 16'hEAFF;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~23_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~22_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~30_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .mask = 16'h3330;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~30 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~30_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~31_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .mask = 16'hAB01;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~31 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .mask = 16'hA2A0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .mask = 16'hB200;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .mask = 16'h5D55;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~5_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .mask = 16'hF0C0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .mask = 16'hEE10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~8_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|I2C_BIT~q ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|comb~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Mux1~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .mask = 16'h32AA;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Mux1~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~7_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~5_combout ),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y10_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X18_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~6_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .mask = 16'h10B0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .mask = 16'hEEFE;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|END~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .mask = 16'h5545;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .mask = 16'h5557;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .mask = 16'h0022;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .mask = 16'h33B3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~3_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .mask = 16'hFEEE;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SCLK~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SDO~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .mask = 16'h8888;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SDO~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .mask = 16'hCBDB;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SDO~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Equal3~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SDO~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .mask = 16'h000D;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|mI2C_WR~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Equal5~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Equal0~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SDO~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SDO~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .mask = 16'hFF02;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|comb~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SDO~3_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SDO~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .mask = 16'hC8CC;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SDO~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X19_Y8_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X19_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X19_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0]~6_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0]~7 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .mask = 16'h33CC;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[0]~7 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X19_Y8_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X19_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X19_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1]~8_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1]~9 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .mask = 16'h3C3F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[1]~9 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X19_Y8_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X19_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X19_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2]~10_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2]~11 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .mask = 16'hC30C;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[2]~11 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X19_Y8_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X19_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X19_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3]~13_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3]~14 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .mask = 16'h3C3F;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[3]~14 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X19_Y8_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X19_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X19_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4]~15_combout ),
	.Cout(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4]~16 ),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .mask = 16'hA50A;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[4]~16 ),
	.Qin(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.Clk(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X19_Y8_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X19_Y8_SIG ),
	.SyncReset(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X19_Y8_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X19_Y8_GND),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~17_combout ),
	.Cout(),
	.Q(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]));
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .mask = 16'h5A5A;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .modeMux = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .BypassEn = 1'b1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SDO~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .mask = 16'h70F0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector2~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .coord_x = 27;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .mask = 16'hBEFF;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector2~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .mask = 16'h8000;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~0_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|END~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .mask = 16'hABAF;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .mask = 16'h0031;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .mask = 16'h05F5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~3_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .mask = 16'hF05C;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .mask = 16'h6084;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SCLK~q ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~5_combout ),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .mask = 16'h5599;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~4_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~6_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector6~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .coord_x = 25;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .mask = 16'hE2CC;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector6~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|Decoder0~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector8~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .mask = 16'hF6FF;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector8~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector9~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .mask = 16'hFDFE;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|Selector9~0_combout ),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|Selector9~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .mask = 16'hFAFA;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|Selector9~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|comb~0 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|comb~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .coord_x = 26;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .mask = 16'h3300;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u0|comb~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u0|comb~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .coord_x = 24;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .mask = 16'hF9CF;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u0|comb~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .mask = 16'h8844;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .mask = 16'h6524;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~1_combout ),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .mask = 16'hCC88;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .mask = 16'h3666;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(vcc),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .mask = 16'h5000;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .mask = 16'h0888;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .mask = 16'hAE10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~6_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .mask = 16'h202A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~7_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~4_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .mask = 16'hFE0E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr0~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .mask = 16'hDE27;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .mask = 16'hF522;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .mask = 16'hF838;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~10_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .mask = 16'h3120;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~11 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .mask = 16'h33C3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .mask = 16'hBF88;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .mask = 16'hB000;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .mask = 16'hB556;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .mask = 16'h6DE2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .mask = 16'hF7FE;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~6_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~7_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .mask = 16'hDD03;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .mask = 16'h8A7C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr10~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .mask = 16'h6106;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .mask = 16'h956A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .mask = 16'hF858;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~10_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .mask = 16'h3120;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~11 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .mask = 16'hE0F8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .mask = 16'hF2F1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~3_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .mask = 16'hE400;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .mask = 16'h9A54;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .mask = 16'h38A8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .mask = 16'h632A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~7_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .mask = 16'hAB89;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .mask = 16'h4010;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr11~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .mask = 16'hBAA0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .mask = 16'hE538;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .mask = 16'h3C80;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .mask = 16'h731A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .mask = 16'h1E4A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .mask = 16'h7F7E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~3_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .mask = 16'hC8D9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .mask = 16'hEA38;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~5_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~6_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .mask = 16'hA2E6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~10_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~7_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .mask = 16'h0A0C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .mask = 16'hB91C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr12~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .mask = 16'h9824;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .mask = 16'h3468;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .mask = 16'h00E4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .mask = 16'h0052;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~2_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .mask = 16'hF4A4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .mask = 16'h54B2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~4_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .mask = 16'h77A0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .mask = 16'hB32C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~6_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .mask = 16'h0081;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .mask = 16'h9102;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~8_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~7_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .mask = 16'hFF80;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr13~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .mask = 16'hD5F6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .mask = 16'h4C42;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .mask = 16'hF6BC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~10_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .mask = 16'hA2E6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .mask = 16'h020A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .mask = 16'h5FFC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~13_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~12_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .mask = 16'h0D01;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .mask = 16'hFFD6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~14_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~15_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .mask = 16'hF0F4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~11_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~16_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .mask = 16'hD9C8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .mask = 16'h3ADE;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .mask = 16'hB6F4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .mask = 16'hFFF2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .mask = 16'h410A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~20_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~19_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .mask = 16'hC2F2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .mask = 16'h8446;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~18_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~22_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~21_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .mask = 16'h3F44;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~17_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~23_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .mask = 16'hEC64;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~24 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~2_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .mask = 16'hF1A1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .mask = 16'h3CB2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~3_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .mask = 16'h1ABA;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .mask = 16'hFAEA;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .mask = 16'h1408;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .mask = 16'h0312;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~8_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~7_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .mask = 16'hBA98;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr14~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .mask = 16'hFF40;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .mask = 16'h0800;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .mask = 16'h3030;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .mask = 16'h8E0E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~3_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .mask = 16'h5F42;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~4_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .mask = 16'h00EC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr1~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .mask = 16'hD35F;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .mask = 16'hEDEC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .mask = 16'h00B8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .mask = 16'h5126;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .mask = 16'hDD11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .mask = 16'hF2A2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .mask = 16'h8B0A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .mask = 16'h94D0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .mask = 16'h9A88;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .mask = 16'h26A6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~5_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~7_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .mask = 16'h38F8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr2~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .mask = 16'h080E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .mask = 16'hF1FE;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .mask = 16'h28FA;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~10_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .mask = 16'hC4E6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~11_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .mask = 16'h00E4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~12 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .mask = 16'h67F6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .mask = 16'hCEC2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .mask = 16'h060C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~4_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .mask = 16'h5FC0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .mask = 16'hE650;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .mask = 16'h0C80;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .mask = 16'h05F8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~7_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .coord_y = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .mask = 16'hA8AD;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr3~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .mask = 16'hFDF8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .mask = 16'hFBDA;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .mask = 16'h00D8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .mask = 16'hAAB1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .mask = 16'h9A80;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .mask = 16'h84A8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .mask = 16'hE6FC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~4_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .mask = 16'hC8CB;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .mask = 16'h61A8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~7_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~3_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .mask = 16'h77A0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~2_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .mask = 16'hBFAA;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr4~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .mask = 16'h5318;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .mask = 16'hBBB8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .mask = 16'hC03F;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .mask = 16'h64E0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~1_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .mask = 16'h9B8A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .mask = 16'hAEEE;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~4_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~3_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .mask = 16'h53F0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .mask = 16'h6E8A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .mask = 16'h70F0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .mask = 16'hCB82;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~7_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .mask = 16'h6F7C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr5~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .mask = 16'h6ECC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .mask = 16'hBE2C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .mask = 16'h5F30;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~10 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~1_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~0_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .mask = 16'h005C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .mask = 16'hF4F2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~3_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .mask = 16'hF0F4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .mask = 16'h1388;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 (
	.A(vcc),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .mask = 16'hC03C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .mask = 16'hB384;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~7_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~6_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .mask = 16'hFC0A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .coord_y = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .mask = 16'hD33E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr6~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .mask = 16'h4C48;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .coord_z = 14;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .mask = 16'h4222;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .mask = 16'h0732;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .mask = 16'hEE05;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(vcc),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .mask = 16'h1100;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~4_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~3_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .mask = 16'h707A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .coord_z = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .mask = 16'h767C;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .mask = 16'hF358;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .coord_z = 4;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .mask = 16'h3FE2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~7_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~8_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .coord_x = 21;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .mask = 16'hA080;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr7~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .mask = 16'h3900;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .mask = 16'h0A28;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .mask = 16'h5804;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .mask = 16'h8A20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .mask = 16'hFE3E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .mask = 16'h46BA;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [0]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~5_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .coord_y = 6;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .coord_z = 15;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .mask = 16'h98DC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .coord_z = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .mask = 16'h0110;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~3_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~7_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .coord_x = 20;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .coord_y = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .coord_z = 1;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .mask = 16'hF588;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr8~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .coord_z = 2;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .mask = 16'h95CA;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~0_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .coord_z = 9;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .mask = 16'h6000;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .coord_z = 0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .mask = 16'h1450;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~1_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~2_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .coord_z = 3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .mask = 16'hCCEC;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~3 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .coord_z = 12;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .mask = 16'hBD7E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .coord_z = 5;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .mask = 16'h9C90;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .coord_z = 10;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .mask = 16'hCF9E;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 (
	.A(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~5_combout ),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [3]),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .coord_z = 13;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .mask = 16'hE0E3;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [6]),
	.B(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [1]),
	.C(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [5]),
	.D(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .coord_z = 8;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .mask = 16'h8478;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 (
	.A(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX [4]),
	.B(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~8_combout ),
	.C(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~4_combout ),
	.D(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~7_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .coord_x = 19;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .coord_y = 7;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .coord_z = 11;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .mask = 16'h770A;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .modeMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .FeedbackMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .ShiftMux = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .BypassEn = 1'b0;
defparam \camera_if_inst|u_I2C_AV_Config|u_I2C_OV7670_Config|WideOr9~9 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|v_cnt[0] (
	.A(\camera_if_inst|v_cnt [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\camera_if_inst|v_cnt [0]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[0]~16_combout ),
	.Cout(\camera_if_inst|v_cnt[0]~17 ),
	.Q(\camera_if_inst|v_cnt [0]));
defparam \camera_if_inst|v_cnt[0] .coord_x = 8;
defparam \camera_if_inst|v_cnt[0] .coord_y = 11;
defparam \camera_if_inst|v_cnt[0] .coord_z = 0;
defparam \camera_if_inst|v_cnt[0] .mask = 16'h55AA;
defparam \camera_if_inst|v_cnt[0] .modeMux = 1'b0;
defparam \camera_if_inst|v_cnt[0] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[0] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[0] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[0] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[10] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [10]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[9]~36 ),
	.Qin(\camera_if_inst|v_cnt [10]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[10]~37_combout ),
	.Cout(\camera_if_inst|v_cnt[10]~38 ),
	.Q(\camera_if_inst|v_cnt [10]));
defparam \camera_if_inst|v_cnt[10] .coord_x = 8;
defparam \camera_if_inst|v_cnt[10] .coord_y = 11;
defparam \camera_if_inst|v_cnt[10] .coord_z = 10;
defparam \camera_if_inst|v_cnt[10] .mask = 16'hC30C;
defparam \camera_if_inst|v_cnt[10] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[10] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[10] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[10] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[10] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[10]~18 (
	.A(\camera_if_inst|Equal3~3_combout ),
	.B(\camera_if_inst|Equal3~4_combout ),
	.C(\camera_if_inst|cam_vsync_r [0]),
	.D(\camera_if_inst|Equal3~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\camera_if_inst|v_cnt[10]~18_combout ),
	.Cout(),
	.Q());
defparam \camera_if_inst|v_cnt[10]~18 .coord_x = 5;
defparam \camera_if_inst|v_cnt[10]~18 .coord_y = 11;
defparam \camera_if_inst|v_cnt[10]~18 .coord_z = 14;
defparam \camera_if_inst|v_cnt[10]~18 .mask = 16'hF0F1;
defparam \camera_if_inst|v_cnt[10]~18 .modeMux = 1'b0;
defparam \camera_if_inst|v_cnt[10]~18 .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[10]~18 .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[10]~18 .BypassEn = 1'b0;
defparam \camera_if_inst|v_cnt[10]~18 .CarryEnb = 1'b1;

alta_slice \camera_if_inst|v_cnt[11] (
	.A(\camera_if_inst|v_cnt [11]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[10]~38 ),
	.Qin(\camera_if_inst|v_cnt [11]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[11]~39_combout ),
	.Cout(\camera_if_inst|v_cnt[11]~40 ),
	.Q(\camera_if_inst|v_cnt [11]));
defparam \camera_if_inst|v_cnt[11] .coord_x = 8;
defparam \camera_if_inst|v_cnt[11] .coord_y = 11;
defparam \camera_if_inst|v_cnt[11] .coord_z = 11;
defparam \camera_if_inst|v_cnt[11] .mask = 16'h5A5F;
defparam \camera_if_inst|v_cnt[11] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[11] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[11] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[11] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[11] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[12] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [12]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[11]~40 ),
	.Qin(\camera_if_inst|v_cnt [12]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[12]~41_combout ),
	.Cout(\camera_if_inst|v_cnt[12]~42 ),
	.Q(\camera_if_inst|v_cnt [12]));
defparam \camera_if_inst|v_cnt[12] .coord_x = 8;
defparam \camera_if_inst|v_cnt[12] .coord_y = 11;
defparam \camera_if_inst|v_cnt[12] .coord_z = 12;
defparam \camera_if_inst|v_cnt[12] .mask = 16'hC30C;
defparam \camera_if_inst|v_cnt[12] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[12] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[12] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[12] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[12] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[13] (
	.A(\camera_if_inst|v_cnt [13]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[12]~42 ),
	.Qin(\camera_if_inst|v_cnt [13]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[13]~43_combout ),
	.Cout(\camera_if_inst|v_cnt[13]~44 ),
	.Q(\camera_if_inst|v_cnt [13]));
defparam \camera_if_inst|v_cnt[13] .coord_x = 8;
defparam \camera_if_inst|v_cnt[13] .coord_y = 11;
defparam \camera_if_inst|v_cnt[13] .coord_z = 13;
defparam \camera_if_inst|v_cnt[13] .mask = 16'h5A5F;
defparam \camera_if_inst|v_cnt[13] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[13] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[13] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[13] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[13] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[14] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [14]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[13]~44 ),
	.Qin(\camera_if_inst|v_cnt [14]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[14]~45_combout ),
	.Cout(\camera_if_inst|v_cnt[14]~46 ),
	.Q(\camera_if_inst|v_cnt [14]));
defparam \camera_if_inst|v_cnt[14] .coord_x = 8;
defparam \camera_if_inst|v_cnt[14] .coord_y = 11;
defparam \camera_if_inst|v_cnt[14] .coord_z = 14;
defparam \camera_if_inst|v_cnt[14] .mask = 16'hC30C;
defparam \camera_if_inst|v_cnt[14] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[14] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[14] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[14] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[14] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[15] (
	.A(\camera_if_inst|v_cnt [15]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[14]~46 ),
	.Qin(\camera_if_inst|v_cnt [15]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[15]~47_combout ),
	.Cout(),
	.Q(\camera_if_inst|v_cnt [15]));
defparam \camera_if_inst|v_cnt[15] .coord_x = 8;
defparam \camera_if_inst|v_cnt[15] .coord_y = 11;
defparam \camera_if_inst|v_cnt[15] .coord_z = 15;
defparam \camera_if_inst|v_cnt[15] .mask = 16'h5A5A;
defparam \camera_if_inst|v_cnt[15] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[15] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[15] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[15] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[15] .CarryEnb = 1'b1;

alta_slice \camera_if_inst|v_cnt[1] (
	.A(\camera_if_inst|v_cnt [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[0]~17 ),
	.Qin(\camera_if_inst|v_cnt [1]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[1]~19_combout ),
	.Cout(\camera_if_inst|v_cnt[1]~20 ),
	.Q(\camera_if_inst|v_cnt [1]));
defparam \camera_if_inst|v_cnt[1] .coord_x = 8;
defparam \camera_if_inst|v_cnt[1] .coord_y = 11;
defparam \camera_if_inst|v_cnt[1] .coord_z = 1;
defparam \camera_if_inst|v_cnt[1] .mask = 16'h5A5F;
defparam \camera_if_inst|v_cnt[1] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[1] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[1] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[1] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[1] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[2] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[1]~20 ),
	.Qin(\camera_if_inst|v_cnt [2]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[2]~21_combout ),
	.Cout(\camera_if_inst|v_cnt[2]~22 ),
	.Q(\camera_if_inst|v_cnt [2]));
defparam \camera_if_inst|v_cnt[2] .coord_x = 8;
defparam \camera_if_inst|v_cnt[2] .coord_y = 11;
defparam \camera_if_inst|v_cnt[2] .coord_z = 2;
defparam \camera_if_inst|v_cnt[2] .mask = 16'hC30C;
defparam \camera_if_inst|v_cnt[2] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[2] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[2] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[2] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[2] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[3] (
	.A(\camera_if_inst|v_cnt [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[2]~22 ),
	.Qin(\camera_if_inst|v_cnt [3]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[3]~23_combout ),
	.Cout(\camera_if_inst|v_cnt[3]~24 ),
	.Q(\camera_if_inst|v_cnt [3]));
defparam \camera_if_inst|v_cnt[3] .coord_x = 8;
defparam \camera_if_inst|v_cnt[3] .coord_y = 11;
defparam \camera_if_inst|v_cnt[3] .coord_z = 3;
defparam \camera_if_inst|v_cnt[3] .mask = 16'h5A5F;
defparam \camera_if_inst|v_cnt[3] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[3] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[3] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[3] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[3] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[4] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[3]~24 ),
	.Qin(\camera_if_inst|v_cnt [4]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[4]~25_combout ),
	.Cout(\camera_if_inst|v_cnt[4]~26 ),
	.Q(\camera_if_inst|v_cnt [4]));
defparam \camera_if_inst|v_cnt[4] .coord_x = 8;
defparam \camera_if_inst|v_cnt[4] .coord_y = 11;
defparam \camera_if_inst|v_cnt[4] .coord_z = 4;
defparam \camera_if_inst|v_cnt[4] .mask = 16'hC30C;
defparam \camera_if_inst|v_cnt[4] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[4] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[4] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[4] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[4] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[5] (
	.A(\camera_if_inst|v_cnt [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[4]~26 ),
	.Qin(\camera_if_inst|v_cnt [5]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[5]~27_combout ),
	.Cout(\camera_if_inst|v_cnt[5]~28 ),
	.Q(\camera_if_inst|v_cnt [5]));
defparam \camera_if_inst|v_cnt[5] .coord_x = 8;
defparam \camera_if_inst|v_cnt[5] .coord_y = 11;
defparam \camera_if_inst|v_cnt[5] .coord_z = 5;
defparam \camera_if_inst|v_cnt[5] .mask = 16'h5A5F;
defparam \camera_if_inst|v_cnt[5] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[5] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[5] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[5] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[5] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[6] (
	.A(\camera_if_inst|v_cnt [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[5]~28 ),
	.Qin(\camera_if_inst|v_cnt [6]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[6]~29_combout ),
	.Cout(\camera_if_inst|v_cnt[6]~30 ),
	.Q(\camera_if_inst|v_cnt [6]));
defparam \camera_if_inst|v_cnt[6] .coord_x = 8;
defparam \camera_if_inst|v_cnt[6] .coord_y = 11;
defparam \camera_if_inst|v_cnt[6] .coord_z = 6;
defparam \camera_if_inst|v_cnt[6] .mask = 16'hA50A;
defparam \camera_if_inst|v_cnt[6] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[6] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[6] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[6] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[6] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[7] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[6]~30 ),
	.Qin(\camera_if_inst|v_cnt [7]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[7]~31_combout ),
	.Cout(\camera_if_inst|v_cnt[7]~32 ),
	.Q(\camera_if_inst|v_cnt [7]));
defparam \camera_if_inst|v_cnt[7] .coord_x = 8;
defparam \camera_if_inst|v_cnt[7] .coord_y = 11;
defparam \camera_if_inst|v_cnt[7] .coord_z = 7;
defparam \camera_if_inst|v_cnt[7] .mask = 16'h3C3F;
defparam \camera_if_inst|v_cnt[7] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[7] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[7] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[7] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[7] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[8] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [8]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[7]~32 ),
	.Qin(\camera_if_inst|v_cnt [8]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[8]~33_combout ),
	.Cout(\camera_if_inst|v_cnt[8]~34 ),
	.Q(\camera_if_inst|v_cnt [8]));
defparam \camera_if_inst|v_cnt[8] .coord_x = 8;
defparam \camera_if_inst|v_cnt[8] .coord_y = 11;
defparam \camera_if_inst|v_cnt[8] .coord_z = 8;
defparam \camera_if_inst|v_cnt[8] .mask = 16'hC30C;
defparam \camera_if_inst|v_cnt[8] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[8] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[8] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[8] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[8] .CarryEnb = 1'b0;

alta_slice \camera_if_inst|v_cnt[9] (
	.A(vcc),
	.B(\camera_if_inst|v_cnt [9]),
	.C(vcc),
	.D(vcc),
	.Cin(\camera_if_inst|v_cnt[8]~34 ),
	.Qin(\camera_if_inst|v_cnt [9]),
	.Clk(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ),
	.AsyncReset(AsyncReset_X5_Y7_GND),
	.SyncReset(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X5_Y7_GND),
	.LutOut(\camera_if_inst|v_cnt[9]~35_combout ),
	.Cout(\camera_if_inst|v_cnt[9]~36 ),
	.Q(\camera_if_inst|v_cnt [9]));
defparam \camera_if_inst|v_cnt[9] .coord_x = 8;
defparam \camera_if_inst|v_cnt[9] .coord_y = 11;
defparam \camera_if_inst|v_cnt[9] .coord_z = 9;
defparam \camera_if_inst|v_cnt[9] .mask = 16'h3C3F;
defparam \camera_if_inst|v_cnt[9] .modeMux = 1'b1;
defparam \camera_if_inst|v_cnt[9] .FeedbackMux = 1'b0;
defparam \camera_if_inst|v_cnt[9] .ShiftMux = 1'b0;
defparam \camera_if_inst|v_cnt[9] .BypassEn = 1'b1;
defparam \camera_if_inst|v_cnt[9] .CarryEnb = 1'b0;

alta_slice clk_25m(
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\clk_25m~q ),
	.Clk(\e_rxclk~input_o_X33_Y16_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\clk_25m~0_combout ),
	.Cout(),
	.Q(\clk_25m~q ));
defparam clk_25m.coord_x = 24;
defparam clk_25m.coord_y = 9;
defparam clk_25m.coord_z = 4;
defparam clk_25m.mask = 16'h0F0F;
defparam clk_25m.modeMux = 1'b0;
defparam clk_25m.FeedbackMux = 1'b1;
defparam clk_25m.ShiftMux = 1'b0;
defparam clk_25m.BypassEn = 1'b0;
defparam clk_25m.CarryEnb = 1'b1;

alta_io_gclk \clk_25m~clkctrl (
	.inclk(\clk_25m~q ),
	.outclk(\clk_25m~clkctrl_outclk ));
defparam \clk_25m~clkctrl .coord_x = 49;
defparam \clk_25m~clkctrl .coord_y = 15;
defparam \clk_25m~clkctrl .coord_z = 4;

alta_clkenctrl clken_ctrl_X10_Y9_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X10_Y9_SIG_VCC ));
defparam clken_ctrl_X10_Y9_N0.coord_x = 16;
defparam clken_ctrl_X10_Y9_N0.coord_y = 13;
defparam clken_ctrl_X10_Y9_N0.coord_z = 0;
defparam clken_ctrl_X10_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X10_Y9_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X10_Y9_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X10_Y9_SIG_VCC ));
defparam clken_ctrl_X10_Y9_N1.coord_x = 16;
defparam clken_ctrl_X10_Y9_N1.coord_y = 13;
defparam clken_ctrl_X10_Y9_N1.coord_z = 1;
defparam clken_ctrl_X10_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X10_Y9_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X11_Y14_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X11_Y14_SIG_VCC ));
defparam clken_ctrl_X11_Y14_N0.coord_x = 9;
defparam clken_ctrl_X11_Y14_N0.coord_y = 14;
defparam clken_ctrl_X11_Y14_N0.coord_z = 0;
defparam clken_ctrl_X11_Y14_N0.ClkMux = 2'b10;
defparam clken_ctrl_X11_Y14_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X11_Y14_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X11_Y14_SIG_SIG ));
defparam clken_ctrl_X11_Y14_N1.coord_x = 9;
defparam clken_ctrl_X11_Y14_N1.coord_y = 14;
defparam clken_ctrl_X11_Y14_N1.coord_z = 1;
defparam clken_ctrl_X11_Y14_N1.ClkMux = 2'b10;
defparam clken_ctrl_X11_Y14_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X11_Y16_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X11_Y16_SIG_VCC ));
defparam clken_ctrl_X11_Y16_N0.coord_x = 16;
defparam clken_ctrl_X11_Y16_N0.coord_y = 15;
defparam clken_ctrl_X11_Y16_N0.coord_z = 0;
defparam clken_ctrl_X11_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X11_Y16_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X11_Y9_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X11_Y9_SIG_VCC ));
defparam clken_ctrl_X11_Y9_N0.coord_x = 16;
defparam clken_ctrl_X11_Y9_N0.coord_y = 12;
defparam clken_ctrl_X11_Y9_N0.coord_z = 0;
defparam clken_ctrl_X11_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X11_Y9_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X11_Y9_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X11_Y9_SIG_VCC ));
defparam clken_ctrl_X11_Y9_N1.coord_x = 16;
defparam clken_ctrl_X11_Y9_N1.coord_y = 12;
defparam clken_ctrl_X11_Y9_N1.coord_z = 1;
defparam clken_ctrl_X11_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X11_Y9_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X12_Y14_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X12_Y14_SIG_VCC ));
defparam clken_ctrl_X12_Y14_N0.coord_x = 10;
defparam clken_ctrl_X12_Y14_N0.coord_y = 14;
defparam clken_ctrl_X12_Y14_N0.coord_z = 0;
defparam clken_ctrl_X12_Y14_N0.ClkMux = 2'b10;
defparam clken_ctrl_X12_Y14_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X12_Y14_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y14_SIG_SIG ));
defparam clken_ctrl_X12_Y14_N1.coord_x = 10;
defparam clken_ctrl_X12_Y14_N1.coord_y = 14;
defparam clken_ctrl_X12_Y14_N1.coord_z = 1;
defparam clken_ctrl_X12_Y14_N1.ClkMux = 2'b10;
defparam clken_ctrl_X12_Y14_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X12_Y16_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X12_Y16_SIG_VCC ));
defparam clken_ctrl_X12_Y16_N0.coord_x = 17;
defparam clken_ctrl_X12_Y16_N0.coord_y = 15;
defparam clken_ctrl_X12_Y16_N0.coord_z = 0;
defparam clken_ctrl_X12_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X12_Y16_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X12_Y18_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X12_Y18_SIG_SIG ));
defparam clken_ctrl_X12_Y18_N0.coord_x = 11;
defparam clken_ctrl_X12_Y18_N0.coord_y = 14;
defparam clken_ctrl_X12_Y18_N0.coord_z = 0;
defparam clken_ctrl_X12_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X12_Y18_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X12_Y18_N1(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X12_Y18_SIG_VCC ));
defparam clken_ctrl_X12_Y18_N1.coord_x = 11;
defparam clken_ctrl_X12_Y18_N1.coord_y = 14;
defparam clken_ctrl_X12_Y18_N1.coord_z = 1;
defparam clken_ctrl_X12_Y18_N1.ClkMux = 2'b10;
defparam clken_ctrl_X12_Y18_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X12_Y9_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ClkOut(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X12_Y9_SIG_SIG ));
defparam clken_ctrl_X12_Y9_N0.coord_x = 15;
defparam clken_ctrl_X12_Y9_N0.coord_y = 11;
defparam clken_ctrl_X12_Y9_N0.coord_z = 0;
defparam clken_ctrl_X12_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X12_Y9_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X12_Y9_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout ),
	.ClkOut(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X12_Y9_SIG_SIG ));
defparam clken_ctrl_X12_Y9_N1.coord_x = 15;
defparam clken_ctrl_X12_Y9_N1.coord_y = 11;
defparam clken_ctrl_X12_Y9_N1.coord_z = 1;
defparam clken_ctrl_X12_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X12_Y9_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X13_Y10_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X13_Y10_SIG_VCC ));
defparam clken_ctrl_X13_Y10_N0.coord_x = 17;
defparam clken_ctrl_X13_Y10_N0.coord_y = 12;
defparam clken_ctrl_X13_Y10_N0.coord_z = 0;
defparam clken_ctrl_X13_Y10_N0.ClkMux = 2'b10;
defparam clken_ctrl_X13_Y10_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X13_Y10_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X13_Y10_SIG_SIG ));
defparam clken_ctrl_X13_Y10_N1.coord_x = 17;
defparam clken_ctrl_X13_Y10_N1.coord_y = 12;
defparam clken_ctrl_X13_Y10_N1.coord_z = 1;
defparam clken_ctrl_X13_Y10_N1.ClkMux = 2'b10;
defparam clken_ctrl_X13_Y10_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X13_Y16_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X13_Y16_SIG_VCC ));
defparam clken_ctrl_X13_Y16_N0.coord_x = 17;
defparam clken_ctrl_X13_Y16_N0.coord_y = 14;
defparam clken_ctrl_X13_Y16_N0.coord_z = 0;
defparam clken_ctrl_X13_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X13_Y16_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X13_Y18_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X13_Y18_SIG_SIG ));
defparam clken_ctrl_X13_Y18_N0.coord_x = 10;
defparam clken_ctrl_X13_Y18_N0.coord_y = 12;
defparam clken_ctrl_X13_Y18_N0.coord_z = 0;
defparam clken_ctrl_X13_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X13_Y18_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X13_Y18_N1(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X13_Y18_SIG_VCC ));
defparam clken_ctrl_X13_Y18_N1.coord_x = 10;
defparam clken_ctrl_X13_Y18_N1.coord_y = 12;
defparam clken_ctrl_X13_Y18_N1.coord_z = 1;
defparam clken_ctrl_X13_Y18_N1.ClkMux = 2'b10;
defparam clken_ctrl_X13_Y18_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X13_Y7_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X13_Y7_SIG_SIG ));
defparam clken_ctrl_X13_Y7_N0.coord_x = 17;
defparam clken_ctrl_X13_Y7_N0.coord_y = 13;
defparam clken_ctrl_X13_Y7_N0.coord_z = 0;
defparam clken_ctrl_X13_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X13_Y7_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X13_Y7_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ClkOut(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X13_Y7_SIG_SIG ));
defparam clken_ctrl_X13_Y7_N1.coord_x = 17;
defparam clken_ctrl_X13_Y7_N1.coord_y = 13;
defparam clken_ctrl_X13_Y7_N1.coord_z = 1;
defparam clken_ctrl_X13_Y7_N1.ClkMux = 2'b10;
defparam clken_ctrl_X13_Y7_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X13_Y9_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout ),
	.ClkOut(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X13_Y9_SIG_SIG ));
defparam clken_ctrl_X13_Y9_N0.coord_x = 16;
defparam clken_ctrl_X13_Y9_N0.coord_y = 11;
defparam clken_ctrl_X13_Y9_N0.coord_z = 0;
defparam clken_ctrl_X13_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X13_Y9_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X13_Y9_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X13_Y9_SIG_VCC ));
defparam clken_ctrl_X13_Y9_N1.coord_x = 16;
defparam clken_ctrl_X13_Y9_N1.coord_y = 11;
defparam clken_ctrl_X13_Y9_N1.coord_z = 1;
defparam clken_ctrl_X13_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X13_Y9_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X14_Y10_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y10_SIG_SIG ));
defparam clken_ctrl_X14_Y10_N0.coord_x = 16;
defparam clken_ctrl_X14_Y10_N0.coord_y = 9;
defparam clken_ctrl_X14_Y10_N0.coord_z = 0;
defparam clken_ctrl_X14_Y10_N0.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y10_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X14_Y10_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X14_Y10_SIG_VCC ));
defparam clken_ctrl_X14_Y10_N1.coord_x = 16;
defparam clken_ctrl_X14_Y10_N1.coord_y = 9;
defparam clken_ctrl_X14_Y10_N1.coord_z = 1;
defparam clken_ctrl_X14_Y10_N1.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y10_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X14_Y11_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X14_Y11_SIG_VCC ));
defparam clken_ctrl_X14_Y11_N0.coord_x = 15;
defparam clken_ctrl_X14_Y11_N0.coord_y = 10;
defparam clken_ctrl_X14_Y11_N0.coord_z = 0;
defparam clken_ctrl_X14_Y11_N0.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y11_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X14_Y14_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X14_Y14_SIG_VCC ));
defparam clken_ctrl_X14_Y14_N0.coord_x = 14;
defparam clken_ctrl_X14_Y14_N0.coord_y = 15;
defparam clken_ctrl_X14_Y14_N0.coord_z = 0;
defparam clken_ctrl_X14_Y14_N0.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y14_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X14_Y16_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X14_Y16_SIG_VCC ));
defparam clken_ctrl_X14_Y16_N0.coord_x = 13;
defparam clken_ctrl_X14_Y16_N0.coord_y = 14;
defparam clken_ctrl_X14_Y16_N0.coord_z = 0;
defparam clken_ctrl_X14_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y16_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X14_Y18_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X14_Y18_SIG_VCC ));
defparam clken_ctrl_X14_Y18_N0.coord_x = 13;
defparam clken_ctrl_X14_Y18_N0.coord_y = 12;
defparam clken_ctrl_X14_Y18_N0.coord_z = 0;
defparam clken_ctrl_X14_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y18_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X14_Y19_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y19_SIG_INV ));
defparam clken_ctrl_X14_Y19_N0.coord_x = 8;
defparam clken_ctrl_X14_Y19_N0.coord_y = 9;
defparam clken_ctrl_X14_Y19_N0.coord_z = 0;
defparam clken_ctrl_X14_Y19_N0.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y19_N0.ClkEnMux = 2'b11;

alta_clkenctrl clken_ctrl_X14_Y20_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_len_reg[10]~35_combout_X14_Y20_SIG_INV ));
defparam clken_ctrl_X14_Y20_N0.coord_x = 8;
defparam clken_ctrl_X14_Y20_N0.coord_y = 10;
defparam clken_ctrl_X14_Y20_N0.coord_z = 0;
defparam clken_ctrl_X14_Y20_N0.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y20_N0.ClkEnMux = 2'b11;

alta_clkenctrl clken_ctrl_X14_Y8_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X14_Y8_SIG_VCC ));
defparam clken_ctrl_X14_Y8_N0.coord_x = 16;
defparam clken_ctrl_X14_Y8_N0.coord_y = 10;
defparam clken_ctrl_X14_Y8_N0.coord_z = 0;
defparam clken_ctrl_X14_Y8_N0.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y8_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X14_Y8_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ));
defparam clken_ctrl_X14_Y8_N1.coord_x = 16;
defparam clken_ctrl_X14_Y8_N1.coord_y = 10;
defparam clken_ctrl_X14_Y8_N1.coord_z = 1;
defparam clken_ctrl_X14_Y8_N1.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y8_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X14_Y9_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ClkOut(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y9_SIG_SIG ));
defparam clken_ctrl_X14_Y9_N0.coord_x = 17;
defparam clken_ctrl_X14_Y9_N0.coord_y = 11;
defparam clken_ctrl_X14_Y9_N0.coord_z = 0;
defparam clken_ctrl_X14_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y9_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X14_Y9_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X14_Y9_SIG_VCC ));
defparam clken_ctrl_X14_Y9_N1.coord_x = 17;
defparam clken_ctrl_X14_Y9_N1.coord_y = 11;
defparam clken_ctrl_X14_Y9_N1.coord_z = 1;
defparam clken_ctrl_X14_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X14_Y9_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X16_Y10_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ));
defparam clken_ctrl_X16_Y10_N0.coord_x = 19;
defparam clken_ctrl_X16_Y10_N0.coord_y = 9;
defparam clken_ctrl_X16_Y10_N0.coord_z = 0;
defparam clken_ctrl_X16_Y10_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y10_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X16_Y11_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|LUT_INDEX[7]~13_combout_X16_Y11_SIG_SIG ));
defparam clken_ctrl_X16_Y11_N0.coord_x = 20;
defparam clken_ctrl_X16_Y11_N0.coord_y = 5;
defparam clken_ctrl_X16_Y11_N0.coord_z = 0;
defparam clken_ctrl_X16_Y11_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y11_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y11_N1(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X16_Y11_SIG_SIG ));
defparam clken_ctrl_X16_Y11_N1.coord_x = 20;
defparam clken_ctrl_X16_Y11_N1.coord_y = 5;
defparam clken_ctrl_X16_Y11_N1.coord_z = 1;
defparam clken_ctrl_X16_Y11_N1.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y11_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y12_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ));
defparam clken_ctrl_X16_Y12_N0.coord_x = 19;
defparam clken_ctrl_X16_Y12_N0.coord_y = 11;
defparam clken_ctrl_X16_Y12_N0.coord_z = 0;
defparam clken_ctrl_X16_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y12_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X16_Y14_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout ),
	.ClkOut(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X16_Y14_SIG_SIG ));
defparam clken_ctrl_X16_Y14_N0.coord_x = 13;
defparam clken_ctrl_X16_Y14_N0.coord_y = 15;
defparam clken_ctrl_X16_Y14_N0.coord_z = 0;
defparam clken_ctrl_X16_Y14_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y14_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y14_N1(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout ),
	.ClkOut(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X16_Y14_SIG_SIG ));
defparam clken_ctrl_X16_Y14_N1.coord_x = 13;
defparam clken_ctrl_X16_Y14_N1.coord_y = 15;
defparam clken_ctrl_X16_Y14_N1.coord_z = 1;
defparam clken_ctrl_X16_Y14_N1.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y14_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y16_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X16_Y16_SIG_VCC ));
defparam clken_ctrl_X16_Y16_N0.coord_x = 15;
defparam clken_ctrl_X16_Y16_N0.coord_y = 15;
defparam clken_ctrl_X16_Y16_N0.coord_z = 0;
defparam clken_ctrl_X16_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y16_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X16_Y16_N1(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X16_Y16_SIG_VCC ));
defparam clken_ctrl_X16_Y16_N1.coord_x = 15;
defparam clken_ctrl_X16_Y16_N1.coord_y = 15;
defparam clken_ctrl_X16_Y16_N1.coord_z = 1;
defparam clken_ctrl_X16_Y16_N1.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y16_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X16_Y17_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena~combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|read_pointer_counter_clk_ena~combout_X16_Y17_SIG_SIG ));
defparam clken_ctrl_X16_Y17_N0.coord_x = 17;
defparam clken_ctrl_X16_Y17_N0.coord_y = 16;
defparam clken_ctrl_X16_Y17_N0.coord_z = 0;
defparam clken_ctrl_X16_Y17_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y17_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y18_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout ),
	.ClkOut(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y18_SIG_SIG ));
defparam clken_ctrl_X16_Y18_N0.coord_x = 14;
defparam clken_ctrl_X16_Y18_N0.coord_y = 14;
defparam clken_ctrl_X16_Y18_N0.coord_z = 0;
defparam clken_ctrl_X16_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y18_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y18_N1(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout ),
	.ClkOut(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y18_SIG_SIG ));
defparam clken_ctrl_X16_Y18_N1.coord_x = 14;
defparam clken_ctrl_X16_Y18_N1.coord_y = 14;
defparam clken_ctrl_X16_Y18_N1.coord_z = 1;
defparam clken_ctrl_X16_Y18_N1.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y18_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y19_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout ),
	.ClkOut(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[1]~0_combout_X16_Y19_SIG_SIG ));
defparam clken_ctrl_X16_Y19_N0.coord_x = 14;
defparam clken_ctrl_X16_Y19_N0.coord_y = 12;
defparam clken_ctrl_X16_Y19_N0.coord_z = 0;
defparam clken_ctrl_X16_Y19_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y19_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y19_N1(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout ),
	.ClkOut(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_ram_gen:attribute_mem_gen:attribute_mem|wdecoder|auto_generated|eq_node[0]~1_combout_X16_Y19_SIG_SIG ));
defparam clken_ctrl_X16_Y19_N1.coord_x = 14;
defparam clken_ctrl_X16_Y19_N1.coord_y = 12;
defparam clken_ctrl_X16_Y19_N1.coord_z = 1;
defparam clken_ctrl_X16_Y19_N1.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y19_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y8_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X16_Y8_SIG_VCC ));
defparam clken_ctrl_X16_Y8_N0.coord_x = 17;
defparam clken_ctrl_X16_Y8_N0.coord_y = 10;
defparam clken_ctrl_X16_Y8_N0.coord_z = 0;
defparam clken_ctrl_X16_Y8_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y8_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X16_Y8_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y8_SIG_SIG ));
defparam clken_ctrl_X16_Y8_N1.coord_x = 17;
defparam clken_ctrl_X16_Y8_N1.coord_y = 10;
defparam clken_ctrl_X16_Y8_N1.coord_z = 1;
defparam clken_ctrl_X16_Y8_N1.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y8_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y9_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ClkOut(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y9_SIG_SIG ));
defparam clken_ctrl_X16_Y9_N0.coord_x = 17;
defparam clken_ctrl_X16_Y9_N0.coord_y = 9;
defparam clken_ctrl_X16_Y9_N0.coord_z = 0;
defparam clken_ctrl_X16_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y9_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X16_Y9_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X16_Y9_SIG_VCC ));
defparam clken_ctrl_X16_Y9_N1.coord_x = 17;
defparam clken_ctrl_X16_Y9_N1.coord_y = 9;
defparam clken_ctrl_X16_Y9_N1.coord_z = 1;
defparam clken_ctrl_X16_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X16_Y9_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y10_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y10_SIG_SIG ));
defparam clken_ctrl_X17_Y10_N0.coord_x = 24;
defparam clken_ctrl_X17_Y10_N0.coord_y = 6;
defparam clken_ctrl_X17_Y10_N0.coord_z = 0;
defparam clken_ctrl_X17_Y10_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y10_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X17_Y11_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X17_Y11_SIG_SIG ));
defparam clken_ctrl_X17_Y11_N0.coord_x = 24;
defparam clken_ctrl_X17_Y11_N0.coord_y = 5;
defparam clken_ctrl_X17_Y11_N0.coord_z = 0;
defparam clken_ctrl_X17_Y11_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y11_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X17_Y11_N1(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X17_Y11_SIG_VCC ));
defparam clken_ctrl_X17_Y11_N1.coord_x = 24;
defparam clken_ctrl_X17_Y11_N1.coord_y = 5;
defparam clken_ctrl_X17_Y11_N1.coord_z = 1;
defparam clken_ctrl_X17_Y11_N1.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y11_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y14_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0_combout ),
	.ClkOut(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|last_buffer_write_address_sig[0]~0_combout_X17_Y14_SIG_SIG ));
defparam clken_ctrl_X17_Y14_N0.coord_x = 12;
defparam clken_ctrl_X17_Y14_N0.coord_y = 15;
defparam clken_ctrl_X17_Y14_N0.coord_z = 0;
defparam clken_ctrl_X17_Y14_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y14_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X17_Y14_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y14_SIG_VCC ));
defparam clken_ctrl_X17_Y14_N1.coord_x = 12;
defparam clken_ctrl_X17_Y14_N1.coord_y = 15;
defparam clken_ctrl_X17_Y14_N1.coord_z = 1;
defparam clken_ctrl_X17_Y14_N1.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y14_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y15_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y15_SIG_VCC ));
defparam clken_ctrl_X17_Y15_N0.coord_x = 5;
defparam clken_ctrl_X17_Y15_N0.coord_y = 15;
defparam clken_ctrl_X17_Y15_N0.coord_z = 0;
defparam clken_ctrl_X17_Y15_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y15_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y15_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17_combout_X17_Y15_SIG_SIG ));
defparam clken_ctrl_X17_Y15_N1.coord_x = 5;
defparam clken_ctrl_X17_Y15_N1.coord_y = 15;
defparam clken_ctrl_X17_Y15_N1.coord_z = 1;
defparam clken_ctrl_X17_Y15_N1.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y15_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X17_Y16_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout_X17_Y16_SIG_SIG ));
defparam clken_ctrl_X17_Y16_N0.coord_x = 7;
defparam clken_ctrl_X17_Y16_N0.coord_y = 17;
defparam clken_ctrl_X17_Y16_N0.coord_z = 0;
defparam clken_ctrl_X17_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y16_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X17_Y17_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X17_Y17_SIG_SIG ));
defparam clken_ctrl_X17_Y17_N0.coord_x = 6;
defparam clken_ctrl_X17_Y17_N0.coord_y = 16;
defparam clken_ctrl_X17_Y17_N0.coord_z = 0;
defparam clken_ctrl_X17_Y17_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y17_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X17_Y17_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y17_SIG_VCC ));
defparam clken_ctrl_X17_Y17_N1.coord_x = 6;
defparam clken_ctrl_X17_Y17_N1.coord_y = 16;
defparam clken_ctrl_X17_Y17_N1.coord_z = 1;
defparam clken_ctrl_X17_Y17_N1.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y17_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y18_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y18_SIG_VCC ));
defparam clken_ctrl_X17_Y18_N0.coord_x = 15;
defparam clken_ctrl_X17_Y18_N0.coord_y = 14;
defparam clken_ctrl_X17_Y18_N0.coord_z = 0;
defparam clken_ctrl_X17_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y18_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y18_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y18_SIG_SIG ));
defparam clken_ctrl_X17_Y18_N1.coord_x = 15;
defparam clken_ctrl_X17_Y18_N1.coord_y = 14;
defparam clken_ctrl_X17_Y18_N1.coord_z = 1;
defparam clken_ctrl_X17_Y18_N1.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y18_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X17_Y19_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y19_SIG_VCC ));
defparam clken_ctrl_X17_Y19_N0.coord_x = 15;
defparam clken_ctrl_X17_Y19_N0.coord_y = 12;
defparam clken_ctrl_X17_Y19_N0.coord_z = 0;
defparam clken_ctrl_X17_Y19_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y19_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y19_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X17_Y19_SIG_SIG ));
defparam clken_ctrl_X17_Y19_N1.coord_x = 15;
defparam clken_ctrl_X17_Y19_N1.coord_y = 12;
defparam clken_ctrl_X17_Y19_N1.coord_z = 1;
defparam clken_ctrl_X17_Y19_N1.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y19_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X17_Y20_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X17_Y20_SIG_VCC ));
defparam clken_ctrl_X17_Y20_N0.coord_x = 14;
defparam clken_ctrl_X17_Y20_N0.coord_y = 16;
defparam clken_ctrl_X17_Y20_N0.coord_z = 0;
defparam clken_ctrl_X17_Y20_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y20_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y9_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X17_Y9_SIG_VCC ));
defparam clken_ctrl_X17_Y9_N0.coord_x = 15;
defparam clken_ctrl_X17_Y9_N0.coord_y = 9;
defparam clken_ctrl_X17_Y9_N0.coord_z = 0;
defparam clken_ctrl_X17_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y9_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X17_Y9_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X17_Y9_SIG_VCC ));
defparam clken_ctrl_X17_Y9_N1.coord_x = 15;
defparam clken_ctrl_X17_Y9_N1.coord_y = 9;
defparam clken_ctrl_X17_Y9_N1.coord_z = 1;
defparam clken_ctrl_X17_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X17_Y9_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X18_Y10_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y10_SIG_SIG ));
defparam clken_ctrl_X18_Y10_N0.coord_x = 25;
defparam clken_ctrl_X18_Y10_N0.coord_y = 6;
defparam clken_ctrl_X18_Y10_N0.coord_z = 0;
defparam clken_ctrl_X18_Y10_N0.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y10_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X18_Y11_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|i2c_negclk~combout_X18_Y11_SIG_SIG ));
defparam clken_ctrl_X18_Y11_N0.coord_x = 25;
defparam clken_ctrl_X18_Y11_N0.coord_y = 5;
defparam clken_ctrl_X18_Y11_N0.coord_z = 0;
defparam clken_ctrl_X18_Y11_N0.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y11_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X18_Y13_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y13_SIG_VCC ));
defparam clken_ctrl_X18_Y13_N0.coord_x = 5;
defparam clken_ctrl_X18_Y13_N0.coord_y = 17;
defparam clken_ctrl_X18_Y13_N0.coord_z = 0;
defparam clken_ctrl_X18_Y13_N0.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y13_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X18_Y13_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout_X18_Y13_SIG_SIG ));
defparam clken_ctrl_X18_Y13_N1.coord_x = 5;
defparam clken_ctrl_X18_Y13_N1.coord_y = 17;
defparam clken_ctrl_X18_Y13_N1.coord_z = 1;
defparam clken_ctrl_X18_Y13_N1.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y13_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X18_Y15_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0]~17_combout_X18_Y15_SIG_SIG ));
defparam clken_ctrl_X18_Y15_N0.coord_x = 6;
defparam clken_ctrl_X18_Y15_N0.coord_y = 15;
defparam clken_ctrl_X18_Y15_N0.coord_z = 0;
defparam clken_ctrl_X18_Y15_N0.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y15_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X18_Y15_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~20_combout_X18_Y15_SIG_SIG ));
defparam clken_ctrl_X18_Y15_N1.coord_x = 6;
defparam clken_ctrl_X18_Y15_N1.coord_y = 15;
defparam clken_ctrl_X18_Y15_N1.coord_z = 1;
defparam clken_ctrl_X18_Y15_N1.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y15_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X18_Y16_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout_X18_Y16_INV_SIG ));
defparam clken_ctrl_X18_Y16_N0.coord_x = 6;
defparam clken_ctrl_X18_Y16_N0.coord_y = 17;
defparam clken_ctrl_X18_Y16_N0.coord_z = 0;
defparam clken_ctrl_X18_Y16_N0.ClkMux = 2'b11;
defparam clken_ctrl_X18_Y16_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X18_Y16_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout_X18_Y16_SIG_SIG ));
defparam clken_ctrl_X18_Y16_N1.coord_x = 6;
defparam clken_ctrl_X18_Y16_N1.coord_y = 17;
defparam clken_ctrl_X18_Y16_N1.coord_z = 1;
defparam clken_ctrl_X18_Y16_N1.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y16_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X18_Y17_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout_X18_Y17_SIG_SIG ));
defparam clken_ctrl_X18_Y17_N0.coord_x = 5;
defparam clken_ctrl_X18_Y17_N0.coord_y = 16;
defparam clken_ctrl_X18_Y17_N0.coord_z = 0;
defparam clken_ctrl_X18_Y17_N0.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y17_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X18_Y17_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~2_combout_X18_Y17_SIG_SIG ));
defparam clken_ctrl_X18_Y17_N1.coord_x = 5;
defparam clken_ctrl_X18_Y17_N1.coord_y = 16;
defparam clken_ctrl_X18_Y17_N1.coord_z = 1;
defparam clken_ctrl_X18_Y17_N1.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y17_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X18_Y18_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X18_Y18_SIG_SIG ));
defparam clken_ctrl_X18_Y18_N0.coord_x = 8;
defparam clken_ctrl_X18_Y18_N0.coord_y = 16;
defparam clken_ctrl_X18_Y18_N0.coord_z = 0;
defparam clken_ctrl_X18_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y18_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X18_Y18_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X18_Y18_SIG_VCC ));
defparam clken_ctrl_X18_Y18_N1.coord_x = 8;
defparam clken_ctrl_X18_Y18_N1.coord_y = 16;
defparam clken_ctrl_X18_Y18_N1.coord_z = 1;
defparam clken_ctrl_X18_Y18_N1.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y18_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X18_Y19_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X18_Y19_SIG_VCC ));
defparam clken_ctrl_X18_Y19_N0.coord_x = 10;
defparam clken_ctrl_X18_Y19_N0.coord_y = 15;
defparam clken_ctrl_X18_Y19_N0.coord_z = 0;
defparam clken_ctrl_X18_Y19_N0.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y19_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X18_Y20_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|Equal2~0_combout_X18_Y20_SIG_SIG ));
defparam clken_ctrl_X18_Y20_N0.coord_x = 13;
defparam clken_ctrl_X18_Y20_N0.coord_y = 16;
defparam clken_ctrl_X18_Y20_N0.coord_z = 0;
defparam clken_ctrl_X18_Y20_N0.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y20_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X18_Y20_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][7]~q_X18_Y20_SIG_SIG ));
defparam clken_ctrl_X18_Y20_N1.coord_x = 13;
defparam clken_ctrl_X18_Y20_N1.coord_y = 16;
defparam clken_ctrl_X18_Y20_N1.coord_z = 1;
defparam clken_ctrl_X18_Y20_N1.ClkMux = 2'b10;
defparam clken_ctrl_X18_Y20_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X19_Y16_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout_X19_Y16_SIG_SIG ));
defparam clken_ctrl_X19_Y16_N0.coord_x = 4;
defparam clken_ctrl_X19_Y16_N0.coord_y = 17;
defparam clken_ctrl_X19_Y16_N0.coord_z = 0;
defparam clken_ctrl_X19_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X19_Y16_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X19_Y16_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout_X19_Y16_SIG_SIG ));
defparam clken_ctrl_X19_Y16_N1.coord_x = 4;
defparam clken_ctrl_X19_Y16_N1.coord_y = 17;
defparam clken_ctrl_X19_Y16_N1.coord_z = 1;
defparam clken_ctrl_X19_Y16_N1.ClkMux = 2'b10;
defparam clken_ctrl_X19_Y16_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X19_Y17_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11]_X19_Y17_SIG_SIG ));
defparam clken_ctrl_X19_Y17_N0.coord_x = 2;
defparam clken_ctrl_X19_Y17_N0.coord_y = 15;
defparam clken_ctrl_X19_Y17_N0.coord_z = 0;
defparam clken_ctrl_X19_Y17_N0.ClkMux = 2'b10;
defparam clken_ctrl_X19_Y17_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X19_Y17_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout_X19_Y17_SIG_SIG ));
defparam clken_ctrl_X19_Y17_N1.coord_x = 2;
defparam clken_ctrl_X19_Y17_N1.coord_y = 15;
defparam clken_ctrl_X19_Y17_N1.coord_z = 1;
defparam clken_ctrl_X19_Y17_N1.ClkMux = 2'b10;
defparam clken_ctrl_X19_Y17_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X19_Y18_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X19_Y18_SIG_SIG ));
defparam clken_ctrl_X19_Y18_N0.coord_x = 7;
defparam clken_ctrl_X19_Y18_N0.coord_y = 15;
defparam clken_ctrl_X19_Y18_N0.coord_z = 0;
defparam clken_ctrl_X19_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X19_Y18_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X19_Y18_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X19_Y18_SIG_INV ));
defparam clken_ctrl_X19_Y18_N1.coord_x = 7;
defparam clken_ctrl_X19_Y18_N1.coord_y = 15;
defparam clken_ctrl_X19_Y18_N1.coord_z = 1;
defparam clken_ctrl_X19_Y18_N1.ClkMux = 2'b10;
defparam clken_ctrl_X19_Y18_N1.ClkEnMux = 2'b11;

alta_clkenctrl clken_ctrl_X19_Y19_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|status_shift_enable~1_combout_X19_Y19_SIG_SIG ));
defparam clken_ctrl_X19_Y19_N0.coord_x = 9;
defparam clken_ctrl_X19_Y19_N0.coord_y = 15;
defparam clken_ctrl_X19_Y19_N0.coord_z = 0;
defparam clken_ctrl_X19_Y19_N0.ClkMux = 2'b10;
defparam clken_ctrl_X19_Y19_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X19_Y8_N1(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(\camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout ),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk__camera_if_inst|u_I2C_AV_Config|u0|SD_COUNTER[5]~12_combout_X19_Y8_SIG_SIG ));
defparam clken_ctrl_X19_Y8_N1.coord_x = 26;
defparam clken_ctrl_X19_Y8_N1.coord_y = 6;
defparam clken_ctrl_X19_Y8_N1.coord_z = 1;
defparam clken_ctrl_X19_Y8_N1.ClkMux = 2'b10;
defparam clken_ctrl_X19_Y8_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X1_Y1_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked ),
	.ClkEn(),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_locked_X1_Y1_SIG_VCC ));
defparam clken_ctrl_X1_Y1_N0.coord_x = 1;
defparam clken_ctrl_X1_Y1_N0.coord_y = 12;
defparam clken_ctrl_X1_Y1_N0.coord_z = 0;
defparam clken_ctrl_X1_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X1_Y1_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X1_Y7_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X1_Y7_SIG_VCC ));
defparam clken_ctrl_X1_Y7_N0.coord_x = 4;
defparam clken_ctrl_X1_Y7_N0.coord_y = 11;
defparam clken_ctrl_X1_Y7_N0.coord_z = 0;
defparam clken_ctrl_X1_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X1_Y7_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X21_Y14_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|always3~4_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ));
defparam clken_ctrl_X21_Y14_N0.coord_x = 21;
defparam clken_ctrl_X21_Y14_N0.coord_y = 12;
defparam clken_ctrl_X21_Y14_N0.coord_z = 0;
defparam clken_ctrl_X21_Y14_N0.ClkMux = 2'b10;
defparam clken_ctrl_X21_Y14_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X21_Y15_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y15_SIG_VCC ));
defparam clken_ctrl_X21_Y15_N0.coord_x = 3;
defparam clken_ctrl_X21_Y15_N0.coord_y = 15;
defparam clken_ctrl_X21_Y15_N0.coord_z = 0;
defparam clken_ctrl_X21_Y15_N0.ClkMux = 2'b10;
defparam clken_ctrl_X21_Y15_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X21_Y16_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q_X21_Y16_SIG_SIG ));
defparam clken_ctrl_X21_Y16_N0.coord_x = 4;
defparam clken_ctrl_X21_Y16_N0.coord_y = 15;
defparam clken_ctrl_X21_Y16_N0.coord_z = 0;
defparam clken_ctrl_X21_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X21_Y16_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X21_Y17_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y17_SIG_VCC ));
defparam clken_ctrl_X21_Y17_N0.coord_x = 1;
defparam clken_ctrl_X21_Y17_N0.coord_y = 15;
defparam clken_ctrl_X21_Y17_N0.coord_z = 0;
defparam clken_ctrl_X21_Y17_N0.ClkMux = 2'b10;
defparam clken_ctrl_X21_Y17_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X21_Y18_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X21_Y18_SIG_VCC ));
defparam clken_ctrl_X21_Y18_N0.coord_x = 9;
defparam clken_ctrl_X21_Y18_N0.coord_y = 16;
defparam clken_ctrl_X21_Y18_N0.coord_z = 0;
defparam clken_ctrl_X21_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X21_Y18_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X21_Y18_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk_X21_Y18_SIG_VCC ));
defparam clken_ctrl_X21_Y18_N1.coord_x = 9;
defparam clken_ctrl_X21_Y18_N1.coord_y = 16;
defparam clken_ctrl_X21_Y18_N1.coord_z = 1;
defparam clken_ctrl_X21_Y18_N1.ClkMux = 2'b10;
defparam clken_ctrl_X21_Y18_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X21_Y19_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X21_Y19_SIG_SIG ));
defparam clken_ctrl_X21_Y19_N0.coord_x = 11;
defparam clken_ctrl_X21_Y19_N0.coord_y = 15;
defparam clken_ctrl_X21_Y19_N0.coord_z = 0;
defparam clken_ctrl_X21_Y19_N0.ClkMux = 2'b10;
defparam clken_ctrl_X21_Y19_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X21_Y20_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X21_Y20_SIG_VCC ));
defparam clken_ctrl_X21_Y20_N0.coord_x = 10;
defparam clken_ctrl_X21_Y20_N0.coord_y = 17;
defparam clken_ctrl_X21_Y20_N0.coord_z = 0;
defparam clken_ctrl_X21_Y20_N0.ClkMux = 2'b10;
defparam clken_ctrl_X21_Y20_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X22_Y14_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|check_sum[8]~47_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y14_SIG_SIG ));
defparam clken_ctrl_X22_Y14_N0.coord_x = 21;
defparam clken_ctrl_X22_Y14_N0.coord_y = 13;
defparam clken_ctrl_X22_Y14_N0.coord_z = 0;
defparam clken_ctrl_X22_Y14_N0.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y14_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X22_Y14_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y14_SIG_SIG ));
defparam clken_ctrl_X22_Y14_N1.coord_x = 21;
defparam clken_ctrl_X22_Y14_N1.coord_y = 13;
defparam clken_ctrl_X22_Y14_N1.coord_z = 1;
defparam clken_ctrl_X22_Y14_N1.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y14_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X22_Y15_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y15_SIG_SIG ));
defparam clken_ctrl_X22_Y15_N0.coord_x = 21;
defparam clken_ctrl_X22_Y15_N0.coord_y = 14;
defparam clken_ctrl_X22_Y15_N0.coord_z = 0;
defparam clken_ctrl_X22_Y15_N0.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y15_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X22_Y15_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|check_sum[8]~47_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y15_SIG_SIG ));
defparam clken_ctrl_X22_Y15_N1.coord_x = 21;
defparam clken_ctrl_X22_Y15_N1.coord_y = 14;
defparam clken_ctrl_X22_Y15_N1.coord_z = 1;
defparam clken_ctrl_X22_Y15_N1.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y15_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X22_Y17_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|WORD_SR[2]~12_combout_X22_Y17_SIG_SIG ));
defparam clken_ctrl_X22_Y17_N0.coord_x = 5;
defparam clken_ctrl_X22_Y17_N0.coord_y = 14;
defparam clken_ctrl_X22_Y17_N0.coord_z = 0;
defparam clken_ctrl_X22_Y17_N0.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y17_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X22_Y17_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|crc_rom_sr|word_counter[3]~10_combout_X22_Y17_SIG_INV ));
defparam clken_ctrl_X22_Y17_N1.coord_x = 5;
defparam clken_ctrl_X22_Y17_N1.coord_y = 14;
defparam clken_ctrl_X22_Y17_N1.coord_z = 1;
defparam clken_ctrl_X22_Y17_N1.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y17_N1.ClkEnMux = 2'b11;

alta_clkenctrl clken_ctrl_X22_Y18_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_val_shift_reg[0]~1_combout_X22_Y18_SIG_SIG ));
defparam clken_ctrl_X22_Y18_N0.coord_x = 8;
defparam clken_ctrl_X22_Y18_N0.coord_y = 15;
defparam clken_ctrl_X22_Y18_N0.coord_z = 0;
defparam clken_ctrl_X22_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y18_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X22_Y18_N1(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|tdo_crc_gen:tdo_crc_calc|lfsr[12]~1_combout_X22_Y18_SIG_INV ));
defparam clken_ctrl_X22_Y18_N1.coord_x = 8;
defparam clken_ctrl_X22_Y18_N1.coord_y = 15;
defparam clken_ctrl_X22_Y18_N1.coord_z = 1;
defparam clken_ctrl_X22_Y18_N1.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y18_N1.ClkEnMux = 2'b11;

alta_clkenctrl clken_ctrl_X22_Y19_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout ),
	.ClkOut(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X22_Y19_SIG_SIG ));
defparam clken_ctrl_X22_Y19_N0.coord_x = 10;
defparam clken_ctrl_X22_Y19_N0.coord_y = 16;
defparam clken_ctrl_X22_Y19_N0.coord_z = 0;
defparam clken_ctrl_X22_Y19_N0.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y19_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X22_Y19_N1(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout ),
	.ClkOut(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X22_Y19_SIG_SIG ));
defparam clken_ctrl_X22_Y19_N1.coord_x = 10;
defparam clken_ctrl_X22_Y19_N1.coord_y = 16;
defparam clken_ctrl_X22_Y19_N1.coord_z = 1;
defparam clken_ctrl_X22_Y19_N1.ClkMux = 2'b10;
defparam clken_ctrl_X22_Y19_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X23_Y16_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y16_SIG_SIG ));
defparam clken_ctrl_X23_Y16_N0.coord_x = 20;
defparam clken_ctrl_X23_Y16_N0.coord_y = 10;
defparam clken_ctrl_X23_Y16_N0.coord_z = 0;
defparam clken_ctrl_X23_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X23_Y16_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X23_Y16_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X23_Y16_SIG_VCC ));
defparam clken_ctrl_X23_Y16_N1.coord_x = 20;
defparam clken_ctrl_X23_Y16_N1.coord_y = 10;
defparam clken_ctrl_X23_Y16_N1.coord_z = 1;
defparam clken_ctrl_X23_Y16_N1.ClkMux = 2'b10;
defparam clken_ctrl_X23_Y16_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X23_Y19_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout ),
	.ClkOut(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|collect_data~combout_X23_Y19_SIG_SIG ));
defparam clken_ctrl_X23_Y19_N0.coord_x = 11;
defparam clken_ctrl_X23_Y19_N0.coord_y = 16;
defparam clken_ctrl_X23_Y19_N0.coord_z = 0;
defparam clken_ctrl_X23_Y19_N0.ClkMux = 2'b10;
defparam clken_ctrl_X23_Y19_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X24_Y12_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X24_Y12_SIG_VCC ));
defparam clken_ctrl_X24_Y12_N0.coord_x = 19;
defparam clken_ctrl_X24_Y12_N0.coord_y = 10;
defparam clken_ctrl_X24_Y12_N0.coord_z = 0;
defparam clken_ctrl_X24_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X24_Y12_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X24_Y15_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|cnt[4]~13_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[4]~13_combout_X24_Y15_SIG_SIG ));
defparam clken_ctrl_X24_Y15_N1.coord_x = 21;
defparam clken_ctrl_X24_Y15_N1.coord_y = 10;
defparam clken_ctrl_X24_Y15_N1.coord_z = 1;
defparam clken_ctrl_X24_Y15_N1.ClkMux = 2'b10;
defparam clken_ctrl_X24_Y15_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X24_Y16_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X24_Y16_SIG_SIG ));
defparam clken_ctrl_X24_Y16_N0.coord_x = 20;
defparam clken_ctrl_X24_Y16_N0.coord_y = 12;
defparam clken_ctrl_X24_Y16_N0.coord_z = 0;
defparam clken_ctrl_X24_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X24_Y16_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X24_Y16_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X24_Y16_SIG_VCC ));
defparam clken_ctrl_X24_Y16_N1.coord_x = 20;
defparam clken_ctrl_X24_Y16_N1.coord_y = 12;
defparam clken_ctrl_X24_Y16_N1.coord_z = 1;
defparam clken_ctrl_X24_Y16_N1.ClkMux = 2'b10;
defparam clken_ctrl_X24_Y16_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X24_Y18_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X24_Y18_SIG_VCC ));
defparam clken_ctrl_X24_Y18_N0.coord_x = 1;
defparam clken_ctrl_X24_Y18_N0.coord_y = 11;
defparam clken_ctrl_X24_Y18_N0.coord_z = 0;
defparam clken_ctrl_X24_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X24_Y18_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X24_Y19_N0(
	.ClkIn(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout ),
	.ClkOut(\altera_internal_jtag~TCKUTAPclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|trigger_setup_ena~combout_X24_Y19_SIG_SIG ));
defparam clken_ctrl_X24_Y19_N0.coord_x = 12;
defparam clken_ctrl_X24_Y19_N0.coord_y = 16;
defparam clken_ctrl_X24_Y19_N0.coord_z = 0;
defparam clken_ctrl_X24_Y19_N0.ClkMux = 2'b10;
defparam clken_ctrl_X24_Y19_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X24_Y19_N1(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout ),
	.ClkOut(\clk~inputclkctrl_outclk__auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|sld_buffer_manager_inst|final_trigger_set~4_combout_X24_Y19_SIG_SIG ));
defparam clken_ctrl_X24_Y19_N1.coord_x = 12;
defparam clken_ctrl_X24_Y19_N1.coord_y = 16;
defparam clken_ctrl_X24_Y19_N1.coord_z = 1;
defparam clken_ctrl_X24_Y19_N1.ClkMux = 2'b10;
defparam clken_ctrl_X24_Y19_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X25_Y12_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|crc32_inst|crc_data[29]~9_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y12_SIG_SIG ));
defparam clken_ctrl_X25_Y12_N0.coord_x = 21;
defparam clken_ctrl_X25_Y12_N0.coord_y = 9;
defparam clken_ctrl_X25_Y12_N0.coord_z = 0;
defparam clken_ctrl_X25_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X25_Y12_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X25_Y12_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X25_Y12_SIG_VCC ));
defparam clken_ctrl_X25_Y12_N1.coord_x = 21;
defparam clken_ctrl_X25_Y12_N1.coord_y = 9;
defparam clken_ctrl_X25_Y12_N1.coord_z = 1;
defparam clken_ctrl_X25_Y12_N1.ClkMux = 2'b10;
defparam clken_ctrl_X25_Y12_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X25_Y13_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|crc32_inst|crc_data[29]~9_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y13_SIG_SIG ));
defparam clken_ctrl_X25_Y13_N0.coord_x = 22;
defparam clken_ctrl_X25_Y13_N0.coord_y = 9;
defparam clken_ctrl_X25_Y13_N0.coord_z = 0;
defparam clken_ctrl_X25_Y13_N0.ClkMux = 2'b10;
defparam clken_ctrl_X25_Y13_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X25_Y13_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout_X25_Y13_SIG_SIG ));
defparam clken_ctrl_X25_Y13_N1.coord_x = 22;
defparam clken_ctrl_X25_Y13_N1.coord_y = 9;
defparam clken_ctrl_X25_Y13_N1.coord_z = 1;
defparam clken_ctrl_X25_Y13_N1.ClkMux = 2'b10;
defparam clken_ctrl_X25_Y13_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X25_Y15_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk_25m~clkctrl_outclk_X25_Y15_SIG_VCC ));
defparam clken_ctrl_X25_Y15_N0.coord_x = 20;
defparam clken_ctrl_X25_Y15_N0.coord_y = 14;
defparam clken_ctrl_X25_Y15_N0.coord_z = 0;
defparam clken_ctrl_X25_Y15_N0.ClkMux = 2'b10;
defparam clken_ctrl_X25_Y15_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X25_Y15_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X25_Y15_SIG_SIG ));
defparam clken_ctrl_X25_Y15_N1.coord_x = 20;
defparam clken_ctrl_X25_Y15_N1.coord_y = 14;
defparam clken_ctrl_X25_Y15_N1.coord_z = 1;
defparam clken_ctrl_X25_Y15_N1.ClkMux = 2'b10;
defparam clken_ctrl_X25_Y15_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X25_Y18_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ));
defparam clken_ctrl_X25_Y18_N0.coord_x = 2;
defparam clken_ctrl_X25_Y18_N0.coord_y = 11;
defparam clken_ctrl_X25_Y18_N0.coord_z = 0;
defparam clken_ctrl_X25_Y18_N0.ClkMux = 2'b10;
defparam clken_ctrl_X25_Y18_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X25_Y19_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ));
defparam clken_ctrl_X25_Y19_N0.coord_x = 2;
defparam clken_ctrl_X25_Y19_N0.coord_y = 12;
defparam clken_ctrl_X25_Y19_N0.coord_z = 0;
defparam clken_ctrl_X25_Y19_N0.ClkMux = 2'b10;
defparam clken_ctrl_X25_Y19_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X26_Y12_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|crc32_inst|crc_data[29]~9_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y12_SIG_SIG ));
defparam clken_ctrl_X26_Y12_N0.coord_x = 20;
defparam clken_ctrl_X26_Y12_N0.coord_y = 9;
defparam clken_ctrl_X26_Y12_N0.coord_z = 0;
defparam clken_ctrl_X26_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X26_Y12_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X26_Y13_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|crc32_inst|crc_data[29]~9_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y13_SIG_SIG ));
defparam clken_ctrl_X26_Y13_N0.coord_x = 22;
defparam clken_ctrl_X26_Y13_N0.coord_y = 8;
defparam clken_ctrl_X26_Y13_N0.coord_z = 0;
defparam clken_ctrl_X26_Y13_N0.ClkMux = 2'b10;
defparam clken_ctrl_X26_Y13_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X26_Y15_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ));
defparam clken_ctrl_X26_Y15_N1.coord_x = 19;
defparam clken_ctrl_X26_Y15_N1.coord_y = 14;
defparam clken_ctrl_X26_Y15_N1.coord_z = 1;
defparam clken_ctrl_X26_Y15_N1.ClkMux = 2'b10;
defparam clken_ctrl_X26_Y15_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X26_Y16_N0(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X26_Y16_SIG_SIG ));
defparam clken_ctrl_X26_Y16_N0.coord_x = 19;
defparam clken_ctrl_X26_Y16_N0.coord_y = 12;
defparam clken_ctrl_X26_Y16_N0.coord_z = 0;
defparam clken_ctrl_X26_Y16_N0.ClkMux = 2'b10;
defparam clken_ctrl_X26_Y16_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X26_Y16_N1(
	.ClkIn(\clk_25m~clkctrl_outclk ),
	.ClkEn(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.ClkOut(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X26_Y16_SIG_SIG ));
defparam clken_ctrl_X26_Y16_N1.coord_x = 19;
defparam clken_ctrl_X26_Y16_N1.coord_y = 12;
defparam clken_ctrl_X26_Y16_N1.coord_z = 1;
defparam clken_ctrl_X26_Y16_N1.ClkMux = 2'b10;
defparam clken_ctrl_X26_Y16_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X28_Y9_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X28_Y9_SIG_VCC ));
defparam clken_ctrl_X28_Y9_N0.coord_x = 24;
defparam clken_ctrl_X28_Y9_N0.coord_y = 8;
defparam clken_ctrl_X28_Y9_N0.coord_z = 0;
defparam clken_ctrl_X28_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X28_Y9_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X29_Y9_N0(
	.ClkIn(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\alt_pll_inst|altpll_component|auto_generated|wire_pll1_clk[0]~clkctrl_outclk_X29_Y9_SIG_VCC ));
defparam clken_ctrl_X29_Y9_N0.coord_x = 25;
defparam clken_ctrl_X29_Y9_N0.coord_y = 8;
defparam clken_ctrl_X29_Y9_N0.coord_z = 0;
defparam clken_ctrl_X29_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X29_Y9_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X2_Y7_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X2_Y7_SIG_VCC ));
defparam clken_ctrl_X2_Y7_N0.coord_x = 5;
defparam clken_ctrl_X2_Y7_N0.coord_y = 11;
defparam clken_ctrl_X2_Y7_N0.coord_z = 0;
defparam clken_ctrl_X2_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X2_Y7_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X33_Y12_N0(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(reset_init[5]),
	.ClkOut(\clk~inputclkctrl_outclk__reset_init[5]_X33_Y12_SIG_INV ));
defparam clken_ctrl_X33_Y12_N0.coord_x = 47;
defparam clken_ctrl_X33_Y12_N0.coord_y = 15;
defparam clken_ctrl_X33_Y12_N0.coord_z = 0;
defparam clken_ctrl_X33_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X33_Y12_N0.ClkEnMux = 2'b11;

alta_clkenctrl clken_ctrl_X33_Y12_N1(
	.ClkIn(\clk~inputclkctrl_outclk ),
	.ClkEn(),
	.ClkOut(\clk~inputclkctrl_outclk_X33_Y12_SIG_VCC ));
defparam clken_ctrl_X33_Y12_N1.coord_x = 47;
defparam clken_ctrl_X33_Y12_N1.coord_y = 15;
defparam clken_ctrl_X33_Y12_N1.coord_z = 1;
defparam clken_ctrl_X33_Y12_N1.ClkMux = 2'b10;
defparam clken_ctrl_X33_Y12_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X33_Y16_N0(
	.ClkIn(\e_rxclk~input_o ),
	.ClkEn(),
	.ClkOut(\e_rxclk~input_o_X33_Y16_INV_VCC ));
defparam clken_ctrl_X33_Y16_N0.coord_x = 24;
defparam clken_ctrl_X33_Y16_N0.coord_y = 9;
defparam clken_ctrl_X33_Y16_N0.coord_z = 0;
defparam clken_ctrl_X33_Y16_N0.ClkMux = 2'b11;
defparam clken_ctrl_X33_Y16_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X33_Y16_N1(
	.ClkIn(\e_rxclk~input_o ),
	.ClkEn(\mii_to_rmii_inst|tx_dv_reg~q ),
	.ClkOut(\e_rxclk~input_o__mii_to_rmii_inst|tx_dv_reg~q_X33_Y16_SIG_SIG ));
defparam clken_ctrl_X33_Y16_N1.coord_x = 24;
defparam clken_ctrl_X33_Y16_N1.coord_y = 9;
defparam clken_ctrl_X33_Y16_N1.coord_z = 1;
defparam clken_ctrl_X33_Y16_N1.ClkMux = 2'b10;
defparam clken_ctrl_X33_Y16_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X5_Y7_N1(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(\camera_if_inst|v_cnt[10]~18_combout ),
	.ClkOut(\cam_pclk~input_o__camera_if_inst|v_cnt[10]~18_combout_X5_Y7_SIG_SIG ));
defparam clken_ctrl_X5_Y7_N1.coord_x = 8;
defparam clken_ctrl_X5_Y7_N1.coord_y = 11;
defparam clken_ctrl_X5_Y7_N1.coord_z = 1;
defparam clken_ctrl_X5_Y7_N1.ClkMux = 2'b10;
defparam clken_ctrl_X5_Y7_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X9_Y7_N0(
	.ClkIn(\cam_pclk~input_o ),
	.ClkEn(),
	.ClkOut(\cam_pclk~input_o_X9_Y7_SIG_VCC ));
defparam clken_ctrl_X9_Y7_N0.coord_x = 10;
defparam clken_ctrl_X9_Y7_N0.coord_y = 11;
defparam clken_ctrl_X9_Y7_N0.coord_z = 0;
defparam clken_ctrl_X9_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X9_Y7_N0.ClkEnMux = 2'b01;

alta_dio \clk~input (
	.padio(clk),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\clk~input_o ),
	.regout());
defparam \clk~input .coord_x = 0;
defparam \clk~input .coord_y = 12;
defparam \clk~input .coord_z = 2;
defparam \clk~input .IN_ASYNC_MODE = 1'b0;
defparam \clk~input .IN_SYNC_MODE = 1'b0;
defparam \clk~input .IN_POWERUP = 1'b0;
defparam \clk~input .IN_ASYNC_DISABLE = 1'b0;
defparam \clk~input .IN_SYNC_DISABLE = 1'b0;
defparam \clk~input .OUT_REG_MODE = 1'b0;
defparam \clk~input .OUT_ASYNC_MODE = 1'b0;
defparam \clk~input .OUT_SYNC_MODE = 1'b0;
defparam \clk~input .OUT_POWERUP = 1'b0;
defparam \clk~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \clk~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \clk~input .OUT_SYNC_DISABLE = 1'b0;
defparam \clk~input .OUT_DDIO = 1'b0;
defparam \clk~input .OE_REG_MODE = 1'b0;
defparam \clk~input .OE_ASYNC_MODE = 1'b0;
defparam \clk~input .OE_SYNC_MODE = 1'b0;
defparam \clk~input .OE_POWERUP = 1'b0;
defparam \clk~input .OE_CLKEN_DISABLE = 1'b0;
defparam \clk~input .OE_ASYNC_DISABLE = 1'b0;
defparam \clk~input .OE_SYNC_DISABLE = 1'b0;
defparam \clk~input .OE_DDIO = 1'b0;
defparam \clk~input .CFG_TRI_INPUT = 1'b0;
defparam \clk~input .CFG_PULL_UP = 1'b0;
defparam \clk~input .CFG_OPEN_DRAIN = 1'b0;
defparam \clk~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \clk~input .CFG_PDRV = 7'b0010000;
defparam \clk~input .CFG_NDRV = 7'b0010000;
defparam \clk~input .CFG_KEEP = 2'b00;
defparam \clk~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \clk~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \clk~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \clk~input .CFG_LVDS_IN_EN = 1'b0;
defparam \clk~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \clk~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \clk~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \clk~input .CFG_OSCDIV = 2'b00;
defparam \clk~input .CFG_ROCTUSR = 1'b0;
defparam \clk~input .CFG_SEL_CUA = 1'b0;
defparam \clk~input .CFG_ROCT_EN = 1'b0;
defparam \clk~input .INPUT_ONLY = 1'b1;
defparam \clk~input .DPCLK_DELAY = 4'b0000;
defparam \clk~input .OUT_DELAY = 1'b0;
defparam \clk~input .IN_DATA_DELAY = 3'b000;
defparam \clk~input .IN_REG_DELAY = 3'b000;

alta_io_gclk \clk~inputclkctrl (
	.inclk(\clk~input_o ),
	.outclk(\clk~inputclkctrl_outclk ));
defparam \clk~inputclkctrl .coord_x = 0;
defparam \clk~inputclkctrl .coord_y = 12;
defparam \clk~inputclkctrl .coord_z = 0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .mask = 16'hAA00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~COUT ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .mask = 16'h0F0F;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [0]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita0~combout ),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita0~COUT ),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .mask = 16'h5555;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[0] .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita0~COUT ),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [1]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~combout ),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~COUT ),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .mask = 16'h3C3F;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit[1] .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [0]),
	.Clk(\cam_pclk~input_o_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [12]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [10]),
	.Clk(\cam_pclk~input_o_X16_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [1]),
	.Clk(\cam_pclk~input_o_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(SyncReset_X14_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y8_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [2]),
	.Clk(\cam_pclk~input_o_X10_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [3]),
	.Clk(\cam_pclk~input_o_X11_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [4]),
	.Clk(\cam_pclk~input_o_X11_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [5]),
	.Clk(\cam_pclk~input_o_X10_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [6]),
	.Clk(\cam_pclk~input_o_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(SyncReset_X17_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X17_Y9_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [7]),
	.Clk(\cam_pclk~input_o_X11_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ),
	.SyncReset(SyncReset_X11_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y9_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [8]),
	.Clk(\cam_pclk~input_o_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(SyncReset_X17_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X17_Y9_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [11]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [9]),
	.Clk(\cam_pclk~input_o_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g[9] .CarryEnb = 1'b1;

alta_bram9k \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 (
	.DataInA({vcc, \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], vcc, \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0], \camera_if_inst|cam_data_r1 [4], \camera_if_inst|cam_data_r1 [0]}),
	.DataInB({1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz}),
	.AddressA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0], vcc}),
	.AddressB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0_combout , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell_combout , vcc, vcc, vcc}),
	.ByteEnA({vcc, vcc}),
	.ByteEnB({1'bz, 1'bz}),
	.DataOutA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutA [0]}),
	.DataOutB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [0]}),
	.Clk0(\cam_pclk~input_o ),
	.ClkEn0(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.AsyncReset0(gnd),
	.Clk1(\clk_25m~clkctrl_outclk ),
	.ClkEn1(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.AsyncReset1(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.WeA(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ReA(gnd),
	.WeB(gnd),
	.ReB(vcc),
	.AddressStallA(gnd),
	.AddressStallB(!\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .coord_x = 18;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .CLKMODE = 2'b10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PACKEDMODE = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_CLKIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_CLKOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_CLKIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_CLKOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_RSTIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_RSTOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_RSTIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_RSTOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_WIDTH = 5'b01110;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_WIDTH = 5'b01000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTA_OUTREG = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .PORTB_OUTREG = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .RSEN_DLY = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .DLYTIME = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0 .INIT_VAL = 9216'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

alta_bram9k \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 (
	.DataInA({vcc, \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [1], \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [1], \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [1], \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [1], vcc, \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [1], \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [1], \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [1], \camera_if_inst|cam_data_r1 [3], \camera_if_inst|cam_data_r1 [1]}),
	.DataInB({1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz}),
	.AddressA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0], vcc}),
	.AddressB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0_combout , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell_combout , vcc, vcc, vcc}),
	.ByteEnA({vcc, vcc}),
	.ByteEnB({1'bz, 1'bz}),
	.DataOutA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutA [0]}),
	.DataOutB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [0]}),
	.Clk0(\cam_pclk~input_o ),
	.ClkEn0(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.AsyncReset0(gnd),
	.Clk1(\clk_25m~clkctrl_outclk ),
	.ClkEn1(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.AsyncReset1(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.WeA(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ReA(gnd),
	.WeB(gnd),
	.ReB(vcc),
	.AddressStallA(gnd),
	.AddressStallB(!\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .coord_x = 18;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .CLKMODE = 2'b10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PACKEDMODE = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_CLKIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_CLKOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_CLKIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_CLKOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_RSTIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_RSTOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_RSTIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_RSTOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_WIDTH = 5'b01110;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_WIDTH = 5'b01000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTA_OUTREG = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .PORTB_OUTREG = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .RSEN_DLY = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .DLYTIME = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1 .INIT_VAL = 9216'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

alta_bram9k \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 (
	.DataInA({vcc, \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [2], \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [2], \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [2], \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [2], vcc, \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [2], \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [2], \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [2], \camera_if_inst|cam_data_r1 [5], \camera_if_inst|cam_data_r1 [2]}),
	.DataInB({1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz}),
	.AddressA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0], vcc}),
	.AddressB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0_combout , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell_combout , vcc, vcc, vcc}),
	.ByteEnA({vcc, vcc}),
	.ByteEnB({1'bz, 1'bz}),
	.DataOutA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutA [0]}),
	.DataOutB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [0]}),
	.Clk0(\cam_pclk~input_o ),
	.ClkEn0(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.AsyncReset0(gnd),
	.Clk1(\clk_25m~clkctrl_outclk ),
	.ClkEn1(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.AsyncReset1(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.WeA(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ReA(gnd),
	.WeB(gnd),
	.ReB(vcc),
	.AddressStallA(gnd),
	.AddressStallB(!\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .coord_x = 18;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .CLKMODE = 2'b10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PACKEDMODE = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_CLKIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_CLKOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_CLKIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_CLKOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_RSTIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_RSTOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_RSTIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_RSTOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_WIDTH = 5'b01110;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_WIDTH = 5'b01000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTA_OUTREG = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .PORTB_OUTREG = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .RSEN_DLY = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .DLYTIME = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2 .INIT_VAL = 9216'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

alta_bram9k \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 (
	.DataInA({vcc, \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [6], vcc, \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [6], \camera_if_inst|cam_data_r1 [7], \camera_if_inst|cam_data_r1 [6]}),
	.DataInB({1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz, 1'bz}),
	.AddressA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0], vcc}),
	.AddressB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0_combout , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q , \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell_combout , vcc, vcc, vcc}),
	.ByteEnA({vcc, vcc}),
	.ByteEnB({1'bz, 1'bz}),
	.DataOutA({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutA [0]}),
	.DataOutB({\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [17], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [16], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [15], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [14], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [13], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [12], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [11], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [10], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [9], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [8], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [7], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [6], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [5], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [4], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [3], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [2], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [1], \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [0]}),
	.Clk0(\cam_pclk~input_o ),
	.ClkEn0(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.AsyncReset0(gnd),
	.Clk1(\clk_25m~clkctrl_outclk ),
	.ClkEn1(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.AsyncReset1(\camera_if_inst|Equal4~0clkctrl_outclk ),
	.WeA(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.ReA(gnd),
	.WeB(gnd),
	.ReB(vcc),
	.AddressStallA(gnd),
	.AddressStallB(!\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .coord_x = 18;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .CLKMODE = 2'b10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PACKEDMODE = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTA_CLKIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTA_CLKOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTB_CLKIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTB_CLKOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTA_RSTIN_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTA_RSTOUT_EN = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTB_RSTIN_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTB_RSTOUT_EN = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTA_WIDTH = 5'b01110;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTB_WIDTH = 5'b01000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTA_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTB_WRITETHRU = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTA_OUTREG = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .PORTB_OUTREG = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .RSEN_DLY = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .DLYTIME = 2'b00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6 .INIT_VAL = 9216'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [0]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1_cout ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .mask = 16'h00DD;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [5]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11_cout ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .mask = 16'h002B;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [6]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [6]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~11_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12_combout ),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~13 ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .mask = 16'h962B;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [7]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14_combout ),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~15 ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .mask = 16'h692B;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [8]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [8]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16_combout ),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~17 ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .mask = 16'h964D;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [9]),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [9]),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .mask = 16'h5AA5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [1]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~1_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3_cout ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .mask = 16'h002B;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [2]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~3_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5_cout ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .mask = 16'h002B;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [3]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~5_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7_cout ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .mask = 16'h004D;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [4]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~7_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9_cout ),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .mask = 16'h002B;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~9 .CarryEnb = 1'b0;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~2_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~3_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~0_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .mask = 16'hFFFE;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~q ),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .mask = 16'h55AA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .mask = 16'h4000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .mask = 16'h1000;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .mask = 16'h0200;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .mask = 16'h0200;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .mask = 16'h0004;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .mask = 16'h0100;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X13_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~1_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .mask = 16'h5A5A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .mask = 16'h00FF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~_wirecell .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ),
	.Clk(\clk_25m~clkctrl_outclk_X13_Y10_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .mask = 16'hF0D2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~q ),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y10_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .mask = 16'hC3F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~2_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.Clk(\clk_25m~clkctrl_outclk_X13_Y10_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .mask = 16'h0FF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ),
	.Clk(\clk_25m~clkctrl_outclk_X13_Y10_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .mask = 16'h3CF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~3_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ),
	.Clk(\clk_25m~clkctrl_outclk_X13_Y10_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .mask = 16'hB4F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~4_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.Clk(\clk_25m~clkctrl_outclk_X13_Y10_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .mask = 16'h0FF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y10_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .mask = 16'h3CF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|cntr_cout[5]~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y10_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .mask = 16'hF078;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~5_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y10_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .mask = 16'h0FF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~6_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~q ),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y10_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .mask = 16'h3CF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [0]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [2]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [1]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X13_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~7_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .mask = 16'h3CC3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|parity6 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [0]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X13_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~10_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .mask = 16'h9669;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [1]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~9_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [2]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|_~8_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .mask = 16'h9966;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|sub_parity7a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a0~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [0]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X13_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .mask = 16'h00FF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a10~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a1~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [1]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X16_Y8_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a2~q ),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X13_Y7_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y7_SIG ),
	.SyncReset(SyncReset_X13_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y7_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a3~q ),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X13_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y10_SIG ),
	.SyncReset(SyncReset_X13_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y10_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a4~q ),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [4]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X13_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y10_SIG ),
	.SyncReset(SyncReset_X13_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X13_Y10_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a5~q ),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a6~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a7~q ),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [7]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ),
	.SyncReset(SyncReset_X14_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y10_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a8~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g1p|counter5a9~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]),
	.Clk(\clk_25m~clkctrl_outclk__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout_X14_Y10_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [0]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor1~combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [0]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor0~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .mask = 16'h33CC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor4~combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [1]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [1]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor1~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor4~combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [2]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor2~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .mask = 16'h9696;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor4~combout ),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [3]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor3~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .mask = 16'h5A5A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [4]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor7~combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [4]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y11_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor4~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor7~combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [5]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y11_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor5~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .mask = 16'hA55A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor7~combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [6]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y11_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor6~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .mask = 16'h55AA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [7]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [7]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y11_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor7~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [8]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y11_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor8~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .mask = 16'hA55A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [9]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y11_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g_gray2bin|xor9~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .mask = 16'h5A5A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_brp|dffe12a[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [0]),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor1~combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [0]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor0~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .mask = 16'h55AA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [2]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor4~combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [1]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [1]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor1~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor4~combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [2]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [2]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor2~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .mask = 16'h9696;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor4~combout ),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [3]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor3~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .mask = 16'h5A5A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [5]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [4]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [6]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor7~combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [4]),
	.Clk(\clk_25m~clkctrl_outclk_X10_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor4~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [5]),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [6]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor7~combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [5]),
	.Clk(\clk_25m~clkctrl_outclk_X10_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor5~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .mask = 16'hA55A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [6]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor7~combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [6]),
	.Clk(\clk_25m~clkctrl_outclk_X10_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor6~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .mask = 16'h0FF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [7]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [8]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [7]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor7~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9]),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [8]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [8]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor8~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .mask = 16'hA55A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9]),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [9]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp_gray2bin|xor9~combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .mask = 16'h55AA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_bwp|dffe12a[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [0]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [0]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(SyncReset_X14_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y8_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [10]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [10]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [1]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [2]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [2]),
	.Clk(\clk_25m~clkctrl_outclk_X10_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [3]),
	.Clk(\clk_25m~clkctrl_outclk_X11_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [4]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [4]),
	.Clk(\clk_25m~clkctrl_outclk_X11_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ),
	.SyncReset(SyncReset_X11_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y9_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [5]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [5]),
	.Clk(\clk_25m~clkctrl_outclk_X10_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ),
	.SyncReset(SyncReset_X10_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X10_Y9_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [6]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [7]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [7]),
	.Clk(\clk_25m~clkctrl_outclk_X11_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [8]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [8]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(SyncReset_X17_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X17_Y9_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|delayed_wrptr_g [9]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [9]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [0]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [0]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [0]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(SyncReset_X14_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y8_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~5_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .mask = 16'h6FF6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [10]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [1]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [1]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [1]),
	.Clk(\clk_25m~clkctrl_outclk_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(SyncReset_X14_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y8_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|data_wire[2]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .mask = 16'h0FF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [5]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [2]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [2]),
	.Clk(\clk_25m~clkctrl_outclk_X10_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ),
	.SyncReset(SyncReset_X10_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X10_Y9_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~3_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .mask = 16'h7DBE;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [3]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3]),
	.Clk(\clk_25m~clkctrl_outclk_X11_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ),
	.SyncReset(SyncReset_X11_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y9_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [4]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [7]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [4]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [7]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [4]),
	.Clk(\clk_25m~clkctrl_outclk_X11_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ),
	.SyncReset(SyncReset_X11_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y9_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~2_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .mask = 16'h7BDE;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [5]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [5]),
	.Clk(\clk_25m~clkctrl_outclk_X10_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ),
	.SyncReset(SyncReset_X10_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X10_Y9_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [6]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [6]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(SyncReset_X17_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X17_Y9_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~1_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .mask = 16'h6FF6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [7]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [7]),
	.Clk(\clk_25m~clkctrl_outclk_X11_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [10]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [8]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [8]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(SyncReset_X17_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X17_Y9_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .mask = 16'h6FF6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe14a [9]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9]),
	.Clk(\clk_25m~clkctrl_outclk_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rs_dgwp|dffpipe13|dffe15a[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~4_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|data_wire[2]~0_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdempty_eq_comp|aneb_result_wire[0]~5_combout ),
	.D(\eth_udp_inst|ip_send_inst|read_data_req~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .mask = 16'hFE00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 (
	.A(\camera_if_inst|cam_hsync_r [1]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|data_wire[2]~0_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .mask = 16'hAAA8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~2_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~1_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .mask = 16'hFFFE;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~4 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .mask = 16'h0400;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .mask = 16'h0100;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .mask = 16'h0100;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .mask = 16'h0400;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .mask = 16'h0200;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_comb_bita1~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5_combout ),
	.Cout(),
	.Q());
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .coord_z = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .mask = 16'h0800;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X12_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~6_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .mask = 16'hA5A5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [10]),
	.Clk(\cam_pclk~input_o_X13_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .mask = 16'hC3F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1]),
	.Clk(\cam_pclk~input_o_X13_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1]~8_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .mask = 16'h78F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.Clk(\cam_pclk~input_o_X13_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2]~7_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .mask = 16'h3CF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~5_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]),
	.Clk(\cam_pclk~input_o_X13_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3]~9_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .mask = 16'hD2F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4]),
	.Clk(\cam_pclk~input_o_X14_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4]~5_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .mask = 16'hD2F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~4_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.Clk(\cam_pclk~input_o_X14_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5]~6_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .mask = 16'h0FF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]),
	.Clk(\cam_pclk~input_o_X13_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6]~3_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .mask = 16'h5AF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~1_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7]),
	.Clk(\cam_pclk~input_o_X13_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7]~4_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .mask = 16'hD2F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~3_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8]),
	.Clk(\cam_pclk~input_o_X13_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8]~1_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .mask = 16'h5A5A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~2_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [9]),
	.Clk(\cam_pclk~input_o_X13_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9]~2_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .mask = 16'h3CF0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2~q ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1~q ),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0~q ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X13_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~7_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .mask = 16'h6699;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|parity8 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0~q ),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X13_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~8_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .mask = 16'h9669;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a0 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1~q ),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X13_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~9_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .mask = 16'h6996;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a1 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [9]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8]),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [10]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2~q ),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|_~0_combout_X13_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|_~10_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2~q ));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .mask = 16'h9966;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|sub_parity9a2 .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .mask = 16'h5555;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [8]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X12_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [12]),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [9]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [11]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(SyncReset_X16_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y9_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ram_address_a [11]),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [11]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .coord_z = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .mask = 16'h5A5A;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[11] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [10]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [12]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [12]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .coord_z = 0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[12] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|cntr_b|counter_reg_bit [1]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [0]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X16_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [1]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [2]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [3]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [4]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .coord_z = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [5]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X14_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y9_SIG ),
	.SyncReset(SyncReset_X14_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y9_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [6]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X12_Y9_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X12_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g1p|counter10a [7]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9]),
	.Clk(\cam_pclk~input_o__cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_wrreq~0_combout_X13_Y7_SIG_SIG ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X13_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [0]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [0]),
	.Clk(\cam_pclk~input_o_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [10]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [10]),
	.Clk(\cam_pclk~input_o_X16_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(SyncReset_X16_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y9_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [1]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [1]),
	.Clk(\cam_pclk~input_o_X14_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [2]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [2]),
	.Clk(\cam_pclk~input_o_X10_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [3]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [3]),
	.Clk(\cam_pclk~input_o_X14_Y8_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .coord_y = 10;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] (
	.A(vcc),
	.B(vcc),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [4]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [4]),
	.Clk(\cam_pclk~input_o_X11_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .mask = 16'hF0F0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [5]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [5]),
	.Clk(\cam_pclk~input_o_X10_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ),
	.SyncReset(SyncReset_X10_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X10_Y9_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [6]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [6]),
	.Clk(\cam_pclk~input_o_X17_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X17_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .coord_x = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .coord_z = 4;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [7]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [7]),
	.Clk(\cam_pclk~input_o_X11_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ),
	.SyncReset(SyncReset_X11_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y9_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] (
	.A(),
	.B(),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [8]),
	.D(),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [8]),
	.Clk(\cam_pclk~input_o_X16_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(SyncReset_X16_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y9_VCC),
	.LutOut(),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .coord_z = 2;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .mask = 16'hFFFF;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .modeMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|rdptr_g [9]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [9]),
	.Clk(\cam_pclk~input_o_X16_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .coord_z = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [3]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [5]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [0]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [2]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [0]),
	.Clk(\cam_pclk~input_o_X14_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y9_SIG ),
	.SyncReset(SyncReset_X14_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y9_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~5_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [0]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .mask = 16'h6FF6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [10]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [10]),
	.Clk(\cam_pclk~input_o_X16_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [10]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .coord_z = 1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [3]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [1]),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [1]),
	.Clk(\cam_pclk~input_o_X14_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y9_SIG ),
	.SyncReset(SyncReset_X14_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X14_Y9_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|data_wire[2]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [1]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .coord_z = 8;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .mask = 16'h3C3C;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [5]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [4]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [2]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [7]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [2]),
	.Clk(\cam_pclk~input_o_X10_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ),
	.SyncReset(SyncReset_X10_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X10_Y9_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~3_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [2]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .coord_z = 14;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .mask = 16'h7DBE;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [3]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [3]),
	.Clk(\cam_pclk~input_o_X14_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X14_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [3]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .coord_y = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .coord_z = 11;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .mask = 16'hFF00;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [7]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [9]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [4]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [6]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [4]),
	.Clk(\cam_pclk~input_o_X11_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ),
	.SyncReset(SyncReset_X11_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X11_Y9_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~2_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [4]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .coord_z = 5;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .mask = 16'h6FF6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [5]),
	.Clk(\cam_pclk~input_o_X10_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X10_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [5]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .coord_y = 13;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .coord_z = 15;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [9]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [11]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [6]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [8]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [6]),
	.Clk(\cam_pclk~input_o_X16_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(SyncReset_X16_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y9_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~1_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [6]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .coord_z = 7;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .mask = 16'h9FF9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [7]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [7]),
	.Clk(\cam_pclk~input_o_X11_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X11_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [7]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .coord_x = 16;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .coord_y = 12;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .mask = 16'hAAAA;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [10]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [10]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [8]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrptr_g [12]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [8]),
	.Clk(\cam_pclk~input_o_X16_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(SyncReset_X16_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X16_Y9_VCC),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|wrfull_eq_comp|aneb_result_wire[0]~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [8]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .coord_z = 6;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .mask = 16'hBE7D;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .FeedbackMux = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .BypassEn = 1'b1;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] (
	.A(vcc),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe18a [9]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [9]),
	.Clk(\cam_pclk~input_o_X16_Y9_SIG_VCC ),
	.AsyncReset(\camera_if_inst|Equal4~0clkctrl_outclk__AsyncReset_X16_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9]~feeder_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a [9]));
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .coord_x = 17;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .coord_y = 9;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .coord_z = 3;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .mask = 16'hCCCC;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|ws_dgrp|dffpipe17|dffe19a[9] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[0] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [9]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [16]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [9]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [0]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y8_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y8_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~14_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [0]));
defparam \cmos1_fifo_inst|q[0] .coord_x = 17;
defparam \cmos1_fifo_inst|q[0] .coord_y = 10;
defparam \cmos1_fifo_inst|q[0] .coord_z = 12;
defparam \cmos1_fifo_inst|q[0] .mask = 16'hD728;
defparam \cmos1_fifo_inst|q[0] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[0] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[0] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[0] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[0] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[10] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [11]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [12]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [11]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [10]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y10_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~4_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [10]));
defparam \cmos1_fifo_inst|q[10] .coord_x = 19;
defparam \cmos1_fifo_inst|q[10] .coord_y = 9;
defparam \cmos1_fifo_inst|q[10] .coord_z = 8;
defparam \cmos1_fifo_inst|q[10] .mask = 16'h9F60;
defparam \cmos1_fifo_inst|q[10] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[10] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[10] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[10] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[10] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[11] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [12]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [12]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [11]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [11]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y10_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~20_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [11]));
defparam \cmos1_fifo_inst|q[11] .coord_x = 19;
defparam \cmos1_fifo_inst|q[11] .coord_y = 9;
defparam \cmos1_fifo_inst|q[11] .coord_z = 12;
defparam \cmos1_fifo_inst|q[11] .mask = 16'hC66C;
defparam \cmos1_fifo_inst|q[11] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[11] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[11] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[11] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[11] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[12] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [12]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [12]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [12]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [12]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y10_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~15_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [12]));
defparam \cmos1_fifo_inst|q[12] .coord_x = 19;
defparam \cmos1_fifo_inst|q[12] .coord_y = 9;
defparam \cmos1_fifo_inst|q[12] .coord_z = 14;
defparam \cmos1_fifo_inst|q[12] .mask = 16'hA66A;
defparam \cmos1_fifo_inst|q[12] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[12] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[12] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[12] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[12] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[13] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [11]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [12]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [12]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [13]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y10_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~31_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [13]));
defparam \cmos1_fifo_inst|q[13] .coord_x = 19;
defparam \cmos1_fifo_inst|q[13] .coord_y = 9;
defparam \cmos1_fifo_inst|q[13] .coord_z = 5;
defparam \cmos1_fifo_inst|q[13] .mask = 16'h96CC;
defparam \cmos1_fifo_inst|q[13] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[13] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[13] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[13] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[13] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[14] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [11]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [12]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [12]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [14]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y10_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~7_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [14]));
defparam \cmos1_fifo_inst|q[14] .coord_x = 19;
defparam \cmos1_fifo_inst|q[14] .coord_y = 9;
defparam \cmos1_fifo_inst|q[14] .coord_z = 10;
defparam \cmos1_fifo_inst|q[14] .mask = 16'h96AA;
defparam \cmos1_fifo_inst|q[14] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[14] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[14] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[14] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[14] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[15] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [13]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [12]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [11]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [15]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~23_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [15]));
defparam \cmos1_fifo_inst|q[15] .coord_x = 19;
defparam \cmos1_fifo_inst|q[15] .coord_y = 11;
defparam \cmos1_fifo_inst|q[15] .coord_z = 10;
defparam \cmos1_fifo_inst|q[15] .mask = 16'h96CC;
defparam \cmos1_fifo_inst|q[15] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[15] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[15] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[15] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[15] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[16] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [13]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [12]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [13]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [16]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~10_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [16]));
defparam \cmos1_fifo_inst|q[16] .coord_x = 19;
defparam \cmos1_fifo_inst|q[16] .coord_y = 11;
defparam \cmos1_fifo_inst|q[16] .coord_z = 3;
defparam \cmos1_fifo_inst|q[16] .mask = 16'h96AA;
defparam \cmos1_fifo_inst|q[16] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[16] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[16] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[16] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[16] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[17] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [13]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [13]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [13]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [17]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~26_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [17]));
defparam \cmos1_fifo_inst|q[17] .coord_x = 19;
defparam \cmos1_fifo_inst|q[17] .coord_y = 11;
defparam \cmos1_fifo_inst|q[17] .coord_z = 6;
defparam \cmos1_fifo_inst|q[17] .mask = 16'h96F0;
defparam \cmos1_fifo_inst|q[17] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[17] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[17] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[17] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[17] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[18] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [14]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [13]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [13]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [18]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~2_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [18]));
defparam \cmos1_fifo_inst|q[18] .coord_x = 19;
defparam \cmos1_fifo_inst|q[18] .coord_y = 11;
defparam \cmos1_fifo_inst|q[18] .coord_z = 13;
defparam \cmos1_fifo_inst|q[18] .mask = 16'h96CC;
defparam \cmos1_fifo_inst|q[18] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[18] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[18] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[18] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[18] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[19] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [14]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [13]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [14]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [19]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~18_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [19]));
defparam \cmos1_fifo_inst|q[19] .coord_x = 19;
defparam \cmos1_fifo_inst|q[19] .coord_y = 11;
defparam \cmos1_fifo_inst|q[19] .coord_z = 12;
defparam \cmos1_fifo_inst|q[19] .mask = 16'h96F0;
defparam \cmos1_fifo_inst|q[19] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[19] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[19] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[19] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[19] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[1] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [9]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [9]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [9]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [1]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y8_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y8_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~30_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [1]));
defparam \cmos1_fifo_inst|q[1] .coord_x = 17;
defparam \cmos1_fifo_inst|q[1] .coord_y = 10;
defparam \cmos1_fifo_inst|q[1] .coord_z = 11;
defparam \cmos1_fifo_inst|q[1] .mask = 16'hC66C;
defparam \cmos1_fifo_inst|q[1] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[1] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[1] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[1] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[1] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[20] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [14]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [14]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [14]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [20]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~9_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [20]));
defparam \cmos1_fifo_inst|q[20] .coord_x = 19;
defparam \cmos1_fifo_inst|q[20] .coord_y = 11;
defparam \cmos1_fifo_inst|q[20] .coord_z = 15;
defparam \cmos1_fifo_inst|q[20] .mask = 16'h96AA;
defparam \cmos1_fifo_inst|q[20] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[20] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[20] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[20] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[20] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[21] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [14]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [13]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [14]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [21]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~24_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [21]));
defparam \cmos1_fifo_inst|q[21] .coord_x = 19;
defparam \cmos1_fifo_inst|q[21] .coord_y = 11;
defparam \cmos1_fifo_inst|q[21] .coord_z = 11;
defparam \cmos1_fifo_inst|q[21] .mask = 16'h96F0;
defparam \cmos1_fifo_inst|q[21] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[21] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[21] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[21] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[21] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[22] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [14]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [13]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [14]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [22]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~0_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [22]));
defparam \cmos1_fifo_inst|q[22] .coord_x = 19;
defparam \cmos1_fifo_inst|q[22] .coord_y = 11;
defparam \cmos1_fifo_inst|q[22] .coord_z = 8;
defparam \cmos1_fifo_inst|q[22] .mask = 16'h96CC;
defparam \cmos1_fifo_inst|q[22] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[22] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[22] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[22] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[22] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[23] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [15]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [13]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [14]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [23]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~16_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [23]));
defparam \cmos1_fifo_inst|q[23] .coord_x = 19;
defparam \cmos1_fifo_inst|q[23] .coord_y = 11;
defparam \cmos1_fifo_inst|q[23] .coord_z = 7;
defparam \cmos1_fifo_inst|q[23] .mask = 16'h9F60;
defparam \cmos1_fifo_inst|q[23] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[23] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[23] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[23] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[23] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[24] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [15]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [15]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [14]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [24]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~8_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [24]));
defparam \cmos1_fifo_inst|q[24] .coord_x = 19;
defparam \cmos1_fifo_inst|q[24] .coord_y = 11;
defparam \cmos1_fifo_inst|q[24] .coord_z = 2;
defparam \cmos1_fifo_inst|q[24] .mask = 16'hB478;
defparam \cmos1_fifo_inst|q[24] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[24] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[24] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[24] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[24] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[25] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [15]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [15]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [15]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [25]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y12_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~25_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [25]));
defparam \cmos1_fifo_inst|q[25] .coord_x = 19;
defparam \cmos1_fifo_inst|q[25] .coord_y = 11;
defparam \cmos1_fifo_inst|q[25] .coord_z = 0;
defparam \cmos1_fifo_inst|q[25] .mask = 16'hA66A;
defparam \cmos1_fifo_inst|q[25] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[25] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[25] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[25] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[25] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[26] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [15]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [15]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [16]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [26]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y8_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y8_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~1_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [26]));
defparam \cmos1_fifo_inst|q[26] .coord_x = 17;
defparam \cmos1_fifo_inst|q[26] .coord_y = 10;
defparam \cmos1_fifo_inst|q[26] .coord_z = 14;
defparam \cmos1_fifo_inst|q[26] .mask = 16'hC66C;
defparam \cmos1_fifo_inst|q[26] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[26] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[26] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[26] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[26] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[27] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [15]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [16]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [16]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [27]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y8_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y8_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~17_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [27]));
defparam \cmos1_fifo_inst|q[27] .coord_x = 17;
defparam \cmos1_fifo_inst|q[27] .coord_y = 10;
defparam \cmos1_fifo_inst|q[27] .coord_z = 13;
defparam \cmos1_fifo_inst|q[27] .mask = 16'hD728;
defparam \cmos1_fifo_inst|q[27] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[27] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[27] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[27] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[27] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[28] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [16]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [16]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [16]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [28]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y8_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y8_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~11_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [28]));
defparam \cmos1_fifo_inst|q[28] .coord_x = 17;
defparam \cmos1_fifo_inst|q[28] .coord_y = 10;
defparam \cmos1_fifo_inst|q[28] .coord_z = 5;
defparam \cmos1_fifo_inst|q[28] .mask = 16'hD278;
defparam \cmos1_fifo_inst|q[28] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[28] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[28] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[28] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[28] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[29] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [16]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [15]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [16]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [29]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y8_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y8_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~27_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [29]));
defparam \cmos1_fifo_inst|q[29] .coord_x = 17;
defparam \cmos1_fifo_inst|q[29] .coord_y = 10;
defparam \cmos1_fifo_inst|q[29] .coord_z = 6;
defparam \cmos1_fifo_inst|q[29] .mask = 16'h9F60;
defparam \cmos1_fifo_inst|q[29] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[29] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[29] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[29] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[29] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[2] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [9]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [9]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [10]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [2]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y8_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y8_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~6_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [2]));
defparam \cmos1_fifo_inst|q[2] .coord_x = 17;
defparam \cmos1_fifo_inst|q[2] .coord_y = 10;
defparam \cmos1_fifo_inst|q[2] .coord_z = 15;
defparam \cmos1_fifo_inst|q[2] .mask = 16'hD278;
defparam \cmos1_fifo_inst|q[2] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[2] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[2] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[2] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[2] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[30] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [16]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [15]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [16]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [30]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y8_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y8_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~3_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [30]));
defparam \cmos1_fifo_inst|q[30] .coord_x = 17;
defparam \cmos1_fifo_inst|q[30] .coord_y = 10;
defparam \cmos1_fifo_inst|q[30] .coord_z = 9;
defparam \cmos1_fifo_inst|q[30] .mask = 16'h9C6C;
defparam \cmos1_fifo_inst|q[30] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[30] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[30] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[30] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[30] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[31] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [15]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [16]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [9]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [31]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y8_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y8_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~19_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [31]));
defparam \cmos1_fifo_inst|q[31] .coord_x = 17;
defparam \cmos1_fifo_inst|q[31] .coord_y = 10;
defparam \cmos1_fifo_inst|q[31] .coord_z = 8;
defparam \cmos1_fifo_inst|q[31] .mask = 16'hD278;
defparam \cmos1_fifo_inst|q[31] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[31] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[31] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[31] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[31] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[3] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [9]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [10]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [10]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [3]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y10_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~22_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [3]));
defparam \cmos1_fifo_inst|q[3] .coord_x = 19;
defparam \cmos1_fifo_inst|q[3] .coord_y = 9;
defparam \cmos1_fifo_inst|q[3] .coord_z = 11;
defparam \cmos1_fifo_inst|q[3] .mask = 16'h96F0;
defparam \cmos1_fifo_inst|q[3] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[3] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[3] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[3] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[3] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[4] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [10]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [10]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [10]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [4]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y10_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~13_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [4]));
defparam \cmos1_fifo_inst|q[4] .coord_x = 19;
defparam \cmos1_fifo_inst|q[4] .coord_y = 9;
defparam \cmos1_fifo_inst|q[4] .coord_z = 7;
defparam \cmos1_fifo_inst|q[4] .mask = 16'h96CC;
defparam \cmos1_fifo_inst|q[4] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[4] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[4] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[4] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[4] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[5] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [10]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [9]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [10]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [5]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y10_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~29_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [5]));
defparam \cmos1_fifo_inst|q[5] .coord_x = 19;
defparam \cmos1_fifo_inst|q[5] .coord_y = 9;
defparam \cmos1_fifo_inst|q[5] .coord_z = 0;
defparam \cmos1_fifo_inst|q[5] .mask = 16'h9A6A;
defparam \cmos1_fifo_inst|q[5] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[5] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[5] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[5] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[5] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[6] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [10]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [10]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [9]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [6]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y10_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~5_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [6]));
defparam \cmos1_fifo_inst|q[6] .coord_x = 19;
defparam \cmos1_fifo_inst|q[6] .coord_y = 9;
defparam \cmos1_fifo_inst|q[6] .coord_z = 2;
defparam \cmos1_fifo_inst|q[6] .mask = 16'h96F0;
defparam \cmos1_fifo_inst|q[6] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[6] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[6] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[6] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[6] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[7] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [9]),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [11]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [10]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [7]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y10_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~21_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [7]));
defparam \cmos1_fifo_inst|q[7] .coord_x = 19;
defparam \cmos1_fifo_inst|q[7] .coord_y = 9;
defparam \cmos1_fifo_inst|q[7] .coord_z = 15;
defparam \cmos1_fifo_inst|q[7] .mask = 16'h96F0;
defparam \cmos1_fifo_inst|q[7] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[7] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[7] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[7] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[7] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[8] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [11]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a6__DataOutB [10]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [11]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [8]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y10_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~12_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [8]));
defparam \cmos1_fifo_inst|q[8] .coord_x = 19;
defparam \cmos1_fifo_inst|q[8] .coord_y = 9;
defparam \cmos1_fifo_inst|q[8] .coord_z = 3;
defparam \cmos1_fifo_inst|q[8] .mask = 16'hC66C;
defparam \cmos1_fifo_inst|q[8] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[8] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[8] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[8] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[8] .CarryEnb = 1'b1;

alta_slice \cmos1_fifo_inst|q[9] (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|valid_rdreq~0_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a2__DataOutB [11]),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a0__DataOutB [11]),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|fifo_ram|ram_block11a1__DataOutB [11]),
	.Cin(),
	.Qin(\cmos1_fifo_inst|q [9]),
	.Clk(\clk_25m~clkctrl_outclk_X16_Y10_SIG_VCC ),
	.AsyncReset(AsyncReset_X16_Y10_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\cmos1_fifo_inst|q~28_combout ),
	.Cout(),
	.Q(\cmos1_fifo_inst|q [9]));
defparam \cmos1_fifo_inst|q[9] .coord_x = 19;
defparam \cmos1_fifo_inst|q[9] .coord_y = 9;
defparam \cmos1_fifo_inst|q[9] .coord_z = 4;
defparam \cmos1_fifo_inst|q[9] .mask = 16'hD728;
defparam \cmos1_fifo_inst|q[9] .modeMux = 1'b0;
defparam \cmos1_fifo_inst|q[9] .FeedbackMux = 1'b0;
defparam \cmos1_fifo_inst|q[9] .ShiftMux = 1'b0;
defparam \cmos1_fifo_inst|q[9] .BypassEn = 1'b0;
defparam \cmos1_fifo_inst|q[9] .CarryEnb = 1'b1;

alta_dio \e_rx[0]~input (
	.padio(e_rx[0]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\e_rx[0]~input_o ),
	.regout());
defparam \e_rx[0]~input .coord_x = 49;
defparam \e_rx[0]~input .coord_y = 19;
defparam \e_rx[0]~input .coord_z = 0;
defparam \e_rx[0]~input .IN_ASYNC_MODE = 1'b0;
defparam \e_rx[0]~input .IN_SYNC_MODE = 1'b0;
defparam \e_rx[0]~input .IN_POWERUP = 1'b0;
defparam \e_rx[0]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \e_rx[0]~input .IN_SYNC_DISABLE = 1'b0;
defparam \e_rx[0]~input .OUT_REG_MODE = 1'b0;
defparam \e_rx[0]~input .OUT_ASYNC_MODE = 1'b0;
defparam \e_rx[0]~input .OUT_SYNC_MODE = 1'b0;
defparam \e_rx[0]~input .OUT_POWERUP = 1'b0;
defparam \e_rx[0]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_rx[0]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_rx[0]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \e_rx[0]~input .OUT_DDIO = 1'b0;
defparam \e_rx[0]~input .OE_REG_MODE = 1'b0;
defparam \e_rx[0]~input .OE_ASYNC_MODE = 1'b0;
defparam \e_rx[0]~input .OE_SYNC_MODE = 1'b0;
defparam \e_rx[0]~input .OE_POWERUP = 1'b0;
defparam \e_rx[0]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \e_rx[0]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \e_rx[0]~input .OE_SYNC_DISABLE = 1'b0;
defparam \e_rx[0]~input .OE_DDIO = 1'b0;
defparam \e_rx[0]~input .CFG_TRI_INPUT = 1'b0;
defparam \e_rx[0]~input .CFG_PULL_UP = 1'b0;
defparam \e_rx[0]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \e_rx[0]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_rx[0]~input .CFG_PDRV = 7'b0011010;
defparam \e_rx[0]~input .CFG_NDRV = 7'b0011000;
defparam \e_rx[0]~input .CFG_KEEP = 2'b00;
defparam \e_rx[0]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_rx[0]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_rx[0]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_rx[0]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \e_rx[0]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_rx[0]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_rx[0]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_rx[0]~input .CFG_OSCDIV = 2'b00;
defparam \e_rx[0]~input .CFG_ROCTUSR = 1'b0;
defparam \e_rx[0]~input .CFG_SEL_CUA = 1'b0;
defparam \e_rx[0]~input .CFG_ROCT_EN = 1'b0;
defparam \e_rx[0]~input .INPUT_ONLY = 1'b0;
defparam \e_rx[0]~input .DPCLK_DELAY = 4'b0000;
defparam \e_rx[0]~input .OUT_DELAY = 1'b0;
defparam \e_rx[0]~input .IN_DATA_DELAY = 3'b000;
defparam \e_rx[0]~input .IN_REG_DELAY = 3'b000;

alta_dio \e_rx[1]~input (
	.padio(e_rx[1]),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\e_rx[1]~input_o ),
	.regout());
defparam \e_rx[1]~input .coord_x = 49;
defparam \e_rx[1]~input .coord_y = 20;
defparam \e_rx[1]~input .coord_z = 2;
defparam \e_rx[1]~input .IN_ASYNC_MODE = 1'b0;
defparam \e_rx[1]~input .IN_SYNC_MODE = 1'b0;
defparam \e_rx[1]~input .IN_POWERUP = 1'b0;
defparam \e_rx[1]~input .IN_ASYNC_DISABLE = 1'b0;
defparam \e_rx[1]~input .IN_SYNC_DISABLE = 1'b0;
defparam \e_rx[1]~input .OUT_REG_MODE = 1'b0;
defparam \e_rx[1]~input .OUT_ASYNC_MODE = 1'b0;
defparam \e_rx[1]~input .OUT_SYNC_MODE = 1'b0;
defparam \e_rx[1]~input .OUT_POWERUP = 1'b0;
defparam \e_rx[1]~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_rx[1]~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_rx[1]~input .OUT_SYNC_DISABLE = 1'b0;
defparam \e_rx[1]~input .OUT_DDIO = 1'b0;
defparam \e_rx[1]~input .OE_REG_MODE = 1'b0;
defparam \e_rx[1]~input .OE_ASYNC_MODE = 1'b0;
defparam \e_rx[1]~input .OE_SYNC_MODE = 1'b0;
defparam \e_rx[1]~input .OE_POWERUP = 1'b0;
defparam \e_rx[1]~input .OE_CLKEN_DISABLE = 1'b0;
defparam \e_rx[1]~input .OE_ASYNC_DISABLE = 1'b0;
defparam \e_rx[1]~input .OE_SYNC_DISABLE = 1'b0;
defparam \e_rx[1]~input .OE_DDIO = 1'b0;
defparam \e_rx[1]~input .CFG_TRI_INPUT = 1'b0;
defparam \e_rx[1]~input .CFG_PULL_UP = 1'b0;
defparam \e_rx[1]~input .CFG_OPEN_DRAIN = 1'b0;
defparam \e_rx[1]~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_rx[1]~input .CFG_PDRV = 7'b0011010;
defparam \e_rx[1]~input .CFG_NDRV = 7'b0011000;
defparam \e_rx[1]~input .CFG_KEEP = 2'b00;
defparam \e_rx[1]~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_rx[1]~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_rx[1]~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_rx[1]~input .CFG_LVDS_IN_EN = 1'b0;
defparam \e_rx[1]~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_rx[1]~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_rx[1]~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_rx[1]~input .CFG_OSCDIV = 2'b00;
defparam \e_rx[1]~input .CFG_ROCTUSR = 1'b0;
defparam \e_rx[1]~input .CFG_SEL_CUA = 1'b0;
defparam \e_rx[1]~input .CFG_ROCT_EN = 1'b0;
defparam \e_rx[1]~input .INPUT_ONLY = 1'b0;
defparam \e_rx[1]~input .DPCLK_DELAY = 4'b0000;
defparam \e_rx[1]~input .OUT_DELAY = 1'b0;
defparam \e_rx[1]~input .IN_DATA_DELAY = 3'b000;
defparam \e_rx[1]~input .IN_REG_DELAY = 3'b000;

alta_dio \e_rxclk~input (
	.padio(e_rxclk),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\e_rxclk~input_o ),
	.regout());
defparam \e_rxclk~input .coord_x = 49;
defparam \e_rxclk~input .coord_y = 27;
defparam \e_rxclk~input .coord_z = 2;
defparam \e_rxclk~input .IN_ASYNC_MODE = 1'b0;
defparam \e_rxclk~input .IN_SYNC_MODE = 1'b0;
defparam \e_rxclk~input .IN_POWERUP = 1'b0;
defparam \e_rxclk~input .IN_ASYNC_DISABLE = 1'b0;
defparam \e_rxclk~input .IN_SYNC_DISABLE = 1'b0;
defparam \e_rxclk~input .OUT_REG_MODE = 1'b0;
defparam \e_rxclk~input .OUT_ASYNC_MODE = 1'b0;
defparam \e_rxclk~input .OUT_SYNC_MODE = 1'b0;
defparam \e_rxclk~input .OUT_POWERUP = 1'b0;
defparam \e_rxclk~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_rxclk~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_rxclk~input .OUT_SYNC_DISABLE = 1'b0;
defparam \e_rxclk~input .OUT_DDIO = 1'b0;
defparam \e_rxclk~input .OE_REG_MODE = 1'b0;
defparam \e_rxclk~input .OE_ASYNC_MODE = 1'b0;
defparam \e_rxclk~input .OE_SYNC_MODE = 1'b0;
defparam \e_rxclk~input .OE_POWERUP = 1'b0;
defparam \e_rxclk~input .OE_CLKEN_DISABLE = 1'b0;
defparam \e_rxclk~input .OE_ASYNC_DISABLE = 1'b0;
defparam \e_rxclk~input .OE_SYNC_DISABLE = 1'b0;
defparam \e_rxclk~input .OE_DDIO = 1'b0;
defparam \e_rxclk~input .CFG_TRI_INPUT = 1'b0;
defparam \e_rxclk~input .CFG_PULL_UP = 1'b0;
defparam \e_rxclk~input .CFG_OPEN_DRAIN = 1'b0;
defparam \e_rxclk~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_rxclk~input .CFG_PDRV = 7'b0011010;
defparam \e_rxclk~input .CFG_NDRV = 7'b0011000;
defparam \e_rxclk~input .CFG_KEEP = 2'b00;
defparam \e_rxclk~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_rxclk~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_rxclk~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_rxclk~input .CFG_LVDS_IN_EN = 1'b0;
defparam \e_rxclk~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_rxclk~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_rxclk~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_rxclk~input .CFG_OSCDIV = 2'b00;
defparam \e_rxclk~input .CFG_ROCTUSR = 1'b0;
defparam \e_rxclk~input .CFG_SEL_CUA = 1'b0;
defparam \e_rxclk~input .CFG_ROCT_EN = 1'b0;
defparam \e_rxclk~input .INPUT_ONLY = 1'b0;
defparam \e_rxclk~input .DPCLK_DELAY = 4'b0000;
defparam \e_rxclk~input .OUT_DELAY = 1'b0;
defparam \e_rxclk~input .IN_DATA_DELAY = 3'b000;
defparam \e_rxclk~input .IN_REG_DELAY = 3'b000;

alta_dio \e_rxdv~input (
	.padio(e_rxdv),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\e_rxdv~input_o ),
	.regout());
defparam \e_rxdv~input .coord_x = 49;
defparam \e_rxdv~input .coord_y = 19;
defparam \e_rxdv~input .coord_z = 3;
defparam \e_rxdv~input .IN_ASYNC_MODE = 1'b0;
defparam \e_rxdv~input .IN_SYNC_MODE = 1'b0;
defparam \e_rxdv~input .IN_POWERUP = 1'b0;
defparam \e_rxdv~input .IN_ASYNC_DISABLE = 1'b0;
defparam \e_rxdv~input .IN_SYNC_DISABLE = 1'b0;
defparam \e_rxdv~input .OUT_REG_MODE = 1'b0;
defparam \e_rxdv~input .OUT_ASYNC_MODE = 1'b0;
defparam \e_rxdv~input .OUT_SYNC_MODE = 1'b0;
defparam \e_rxdv~input .OUT_POWERUP = 1'b0;
defparam \e_rxdv~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_rxdv~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_rxdv~input .OUT_SYNC_DISABLE = 1'b0;
defparam \e_rxdv~input .OUT_DDIO = 1'b0;
defparam \e_rxdv~input .OE_REG_MODE = 1'b0;
defparam \e_rxdv~input .OE_ASYNC_MODE = 1'b0;
defparam \e_rxdv~input .OE_SYNC_MODE = 1'b0;
defparam \e_rxdv~input .OE_POWERUP = 1'b0;
defparam \e_rxdv~input .OE_CLKEN_DISABLE = 1'b0;
defparam \e_rxdv~input .OE_ASYNC_DISABLE = 1'b0;
defparam \e_rxdv~input .OE_SYNC_DISABLE = 1'b0;
defparam \e_rxdv~input .OE_DDIO = 1'b0;
defparam \e_rxdv~input .CFG_TRI_INPUT = 1'b0;
defparam \e_rxdv~input .CFG_PULL_UP = 1'b0;
defparam \e_rxdv~input .CFG_OPEN_DRAIN = 1'b0;
defparam \e_rxdv~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_rxdv~input .CFG_PDRV = 7'b0011010;
defparam \e_rxdv~input .CFG_NDRV = 7'b0011000;
defparam \e_rxdv~input .CFG_KEEP = 2'b00;
defparam \e_rxdv~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_rxdv~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_rxdv~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_rxdv~input .CFG_LVDS_IN_EN = 1'b0;
defparam \e_rxdv~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_rxdv~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_rxdv~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_rxdv~input .CFG_OSCDIV = 2'b00;
defparam \e_rxdv~input .CFG_ROCTUSR = 1'b0;
defparam \e_rxdv~input .CFG_SEL_CUA = 1'b0;
defparam \e_rxdv~input .CFG_ROCT_EN = 1'b0;
defparam \e_rxdv~input .INPUT_ONLY = 1'b0;
defparam \e_rxdv~input .DPCLK_DELAY = 4'b0000;
defparam \e_rxdv~input .OUT_DELAY = 1'b0;
defparam \e_rxdv~input .IN_DATA_DELAY = 3'b000;
defparam \e_rxdv~input .IN_REG_DELAY = 3'b000;

alta_dio \e_rxer~input (
	.padio(e_rxer),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\e_rxer~input_o ),
	.regout());
defparam \e_rxer~input .coord_x = 49;
defparam \e_rxer~input .coord_y = 19;
defparam \e_rxer~input .coord_z = 1;
defparam \e_rxer~input .IN_ASYNC_MODE = 1'b0;
defparam \e_rxer~input .IN_SYNC_MODE = 1'b0;
defparam \e_rxer~input .IN_POWERUP = 1'b0;
defparam \e_rxer~input .IN_ASYNC_DISABLE = 1'b0;
defparam \e_rxer~input .IN_SYNC_DISABLE = 1'b0;
defparam \e_rxer~input .OUT_REG_MODE = 1'b0;
defparam \e_rxer~input .OUT_ASYNC_MODE = 1'b0;
defparam \e_rxer~input .OUT_SYNC_MODE = 1'b0;
defparam \e_rxer~input .OUT_POWERUP = 1'b0;
defparam \e_rxer~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_rxer~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_rxer~input .OUT_SYNC_DISABLE = 1'b0;
defparam \e_rxer~input .OUT_DDIO = 1'b0;
defparam \e_rxer~input .OE_REG_MODE = 1'b0;
defparam \e_rxer~input .OE_ASYNC_MODE = 1'b0;
defparam \e_rxer~input .OE_SYNC_MODE = 1'b0;
defparam \e_rxer~input .OE_POWERUP = 1'b0;
defparam \e_rxer~input .OE_CLKEN_DISABLE = 1'b0;
defparam \e_rxer~input .OE_ASYNC_DISABLE = 1'b0;
defparam \e_rxer~input .OE_SYNC_DISABLE = 1'b0;
defparam \e_rxer~input .OE_DDIO = 1'b0;
defparam \e_rxer~input .CFG_TRI_INPUT = 1'b0;
defparam \e_rxer~input .CFG_PULL_UP = 1'b0;
defparam \e_rxer~input .CFG_OPEN_DRAIN = 1'b0;
defparam \e_rxer~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_rxer~input .CFG_PDRV = 7'b0011010;
defparam \e_rxer~input .CFG_NDRV = 7'b0011000;
defparam \e_rxer~input .CFG_KEEP = 2'b00;
defparam \e_rxer~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_rxer~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_rxer~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_rxer~input .CFG_LVDS_IN_EN = 1'b0;
defparam \e_rxer~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_rxer~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_rxer~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_rxer~input .CFG_OSCDIV = 2'b00;
defparam \e_rxer~input .CFG_ROCTUSR = 1'b0;
defparam \e_rxer~input .CFG_SEL_CUA = 1'b0;
defparam \e_rxer~input .CFG_ROCT_EN = 1'b0;
defparam \e_rxer~input .INPUT_ONLY = 1'b0;
defparam \e_rxer~input .DPCLK_DELAY = 4'b0000;
defparam \e_rxer~input .OUT_DELAY = 1'b0;
defparam \e_rxer~input .IN_DATA_DELAY = 3'b000;
defparam \e_rxer~input .IN_REG_DELAY = 3'b000;

alta_dio \e_tx[0]~output (
	.padio(e_tx[0]),
	.datain(\mii_to_rmii_inst|eth_tx_data [0]),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \e_tx[0]~output .coord_x = 49;
defparam \e_tx[0]~output .coord_y = 27;
defparam \e_tx[0]~output .coord_z = 1;
defparam \e_tx[0]~output .IN_ASYNC_MODE = 1'b0;
defparam \e_tx[0]~output .IN_SYNC_MODE = 1'b0;
defparam \e_tx[0]~output .IN_POWERUP = 1'b0;
defparam \e_tx[0]~output .IN_ASYNC_DISABLE = 1'b0;
defparam \e_tx[0]~output .IN_SYNC_DISABLE = 1'b0;
defparam \e_tx[0]~output .OUT_REG_MODE = 1'b0;
defparam \e_tx[0]~output .OUT_ASYNC_MODE = 1'b0;
defparam \e_tx[0]~output .OUT_SYNC_MODE = 1'b0;
defparam \e_tx[0]~output .OUT_POWERUP = 1'b0;
defparam \e_tx[0]~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_tx[0]~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_tx[0]~output .OUT_SYNC_DISABLE = 1'b0;
defparam \e_tx[0]~output .OUT_DDIO = 1'b0;
defparam \e_tx[0]~output .OE_REG_MODE = 1'b0;
defparam \e_tx[0]~output .OE_ASYNC_MODE = 1'b0;
defparam \e_tx[0]~output .OE_SYNC_MODE = 1'b0;
defparam \e_tx[0]~output .OE_POWERUP = 1'b0;
defparam \e_tx[0]~output .OE_CLKEN_DISABLE = 1'b0;
defparam \e_tx[0]~output .OE_ASYNC_DISABLE = 1'b0;
defparam \e_tx[0]~output .OE_SYNC_DISABLE = 1'b0;
defparam \e_tx[0]~output .OE_DDIO = 1'b0;
defparam \e_tx[0]~output .CFG_TRI_INPUT = 1'b0;
defparam \e_tx[0]~output .CFG_PULL_UP = 1'b0;
defparam \e_tx[0]~output .CFG_OPEN_DRAIN = 1'b0;
defparam \e_tx[0]~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_tx[0]~output .CFG_PDRV = 7'b0011010;
defparam \e_tx[0]~output .CFG_NDRV = 7'b0011000;
defparam \e_tx[0]~output .CFG_KEEP = 2'b00;
defparam \e_tx[0]~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_tx[0]~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_tx[0]~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_tx[0]~output .CFG_LVDS_IN_EN = 1'b0;
defparam \e_tx[0]~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_tx[0]~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_tx[0]~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_tx[0]~output .CFG_OSCDIV = 2'b00;
defparam \e_tx[0]~output .CFG_ROCTUSR = 1'b0;
defparam \e_tx[0]~output .CFG_SEL_CUA = 1'b0;
defparam \e_tx[0]~output .CFG_ROCT_EN = 1'b0;
defparam \e_tx[0]~output .INPUT_ONLY = 1'b0;
defparam \e_tx[0]~output .DPCLK_DELAY = 4'b0000;
defparam \e_tx[0]~output .OUT_DELAY = 1'b0;
defparam \e_tx[0]~output .IN_DATA_DELAY = 3'b000;
defparam \e_tx[0]~output .IN_REG_DELAY = 3'b000;

alta_dio \e_tx[1]~output (
	.padio(e_tx[1]),
	.datain(\mii_to_rmii_inst|eth_tx_data [1]),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \e_tx[1]~output .coord_x = 44;
defparam \e_tx[1]~output .coord_y = 29;
defparam \e_tx[1]~output .coord_z = 2;
defparam \e_tx[1]~output .IN_ASYNC_MODE = 1'b0;
defparam \e_tx[1]~output .IN_SYNC_MODE = 1'b0;
defparam \e_tx[1]~output .IN_POWERUP = 1'b0;
defparam \e_tx[1]~output .IN_ASYNC_DISABLE = 1'b0;
defparam \e_tx[1]~output .IN_SYNC_DISABLE = 1'b0;
defparam \e_tx[1]~output .OUT_REG_MODE = 1'b0;
defparam \e_tx[1]~output .OUT_ASYNC_MODE = 1'b0;
defparam \e_tx[1]~output .OUT_SYNC_MODE = 1'b0;
defparam \e_tx[1]~output .OUT_POWERUP = 1'b0;
defparam \e_tx[1]~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_tx[1]~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_tx[1]~output .OUT_SYNC_DISABLE = 1'b0;
defparam \e_tx[1]~output .OUT_DDIO = 1'b0;
defparam \e_tx[1]~output .OE_REG_MODE = 1'b0;
defparam \e_tx[1]~output .OE_ASYNC_MODE = 1'b0;
defparam \e_tx[1]~output .OE_SYNC_MODE = 1'b0;
defparam \e_tx[1]~output .OE_POWERUP = 1'b0;
defparam \e_tx[1]~output .OE_CLKEN_DISABLE = 1'b0;
defparam \e_tx[1]~output .OE_ASYNC_DISABLE = 1'b0;
defparam \e_tx[1]~output .OE_SYNC_DISABLE = 1'b0;
defparam \e_tx[1]~output .OE_DDIO = 1'b0;
defparam \e_tx[1]~output .CFG_TRI_INPUT = 1'b0;
defparam \e_tx[1]~output .CFG_PULL_UP = 1'b0;
defparam \e_tx[1]~output .CFG_OPEN_DRAIN = 1'b0;
defparam \e_tx[1]~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_tx[1]~output .CFG_PDRV = 7'b0011010;
defparam \e_tx[1]~output .CFG_NDRV = 7'b0011000;
defparam \e_tx[1]~output .CFG_KEEP = 2'b00;
defparam \e_tx[1]~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_tx[1]~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_tx[1]~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_tx[1]~output .CFG_LVDS_IN_EN = 1'b0;
defparam \e_tx[1]~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_tx[1]~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_tx[1]~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_tx[1]~output .CFG_OSCDIV = 2'b00;
defparam \e_tx[1]~output .CFG_ROCTUSR = 1'b0;
defparam \e_tx[1]~output .CFG_SEL_CUA = 1'b0;
defparam \e_tx[1]~output .CFG_ROCT_EN = 1'b0;
defparam \e_tx[1]~output .INPUT_ONLY = 1'b0;
defparam \e_tx[1]~output .DPCLK_DELAY = 4'b0000;
defparam \e_tx[1]~output .OUT_DELAY = 1'b0;
defparam \e_tx[1]~output .IN_DATA_DELAY = 3'b000;
defparam \e_tx[1]~output .IN_REG_DELAY = 3'b000;

alta_dio \e_txen~output (
	.padio(e_txen),
	.datain(\mii_to_rmii_inst|eth_tx_dv~q ),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \e_txen~output .coord_x = 43;
defparam \e_txen~output .coord_y = 29;
defparam \e_txen~output .coord_z = 1;
defparam \e_txen~output .IN_ASYNC_MODE = 1'b0;
defparam \e_txen~output .IN_SYNC_MODE = 1'b0;
defparam \e_txen~output .IN_POWERUP = 1'b0;
defparam \e_txen~output .IN_ASYNC_DISABLE = 1'b0;
defparam \e_txen~output .IN_SYNC_DISABLE = 1'b0;
defparam \e_txen~output .OUT_REG_MODE = 1'b0;
defparam \e_txen~output .OUT_ASYNC_MODE = 1'b0;
defparam \e_txen~output .OUT_SYNC_MODE = 1'b0;
defparam \e_txen~output .OUT_POWERUP = 1'b0;
defparam \e_txen~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \e_txen~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \e_txen~output .OUT_SYNC_DISABLE = 1'b0;
defparam \e_txen~output .OUT_DDIO = 1'b0;
defparam \e_txen~output .OE_REG_MODE = 1'b0;
defparam \e_txen~output .OE_ASYNC_MODE = 1'b0;
defparam \e_txen~output .OE_SYNC_MODE = 1'b0;
defparam \e_txen~output .OE_POWERUP = 1'b0;
defparam \e_txen~output .OE_CLKEN_DISABLE = 1'b0;
defparam \e_txen~output .OE_ASYNC_DISABLE = 1'b0;
defparam \e_txen~output .OE_SYNC_DISABLE = 1'b0;
defparam \e_txen~output .OE_DDIO = 1'b0;
defparam \e_txen~output .CFG_TRI_INPUT = 1'b0;
defparam \e_txen~output .CFG_PULL_UP = 1'b0;
defparam \e_txen~output .CFG_OPEN_DRAIN = 1'b0;
defparam \e_txen~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \e_txen~output .CFG_PDRV = 7'b0011010;
defparam \e_txen~output .CFG_NDRV = 7'b0011000;
defparam \e_txen~output .CFG_KEEP = 2'b00;
defparam \e_txen~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \e_txen~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \e_txen~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \e_txen~output .CFG_LVDS_IN_EN = 1'b0;
defparam \e_txen~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \e_txen~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \e_txen~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \e_txen~output .CFG_OSCDIV = 2'b00;
defparam \e_txen~output .CFG_ROCTUSR = 1'b0;
defparam \e_txen~output .CFG_SEL_CUA = 1'b0;
defparam \e_txen~output .CFG_ROCT_EN = 1'b0;
defparam \e_txen~output .INPUT_ONLY = 1'b0;
defparam \e_txen~output .DPCLK_DELAY = 4'b0000;
defparam \e_txen~output .OUT_DELAY = 1'b0;
defparam \e_txen~output .IN_DATA_DELAY = 3'b000;
defparam \e_txen~output .IN_REG_DELAY = 3'b000;

alta_slice \eth_udp_inst|crc32_inst|crc_data[0] (
	.A(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.B(vcc),
	.C(\eth_udp_inst|crc32_inst|crc_data [28]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [0]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~25_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [0]));
defparam \eth_udp_inst|crc32_inst|crc_data[0] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .coord_y = 8;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .coord_z = 14;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .mask = 16'h0550;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[0] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[10] (
	.A(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.B(\eth_udp_inst|crc32_inst|crc_data [6]),
	.C(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.D(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [10]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~30_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [10]));
defparam \eth_udp_inst|crc32_inst|crc_data[10] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .coord_y = 8;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .coord_z = 3;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .mask = 16'h0609;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[10] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[11] (
	.A(\eth_udp_inst|crc32_inst|crc_data [7]),
	.B(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.C(vcc),
	.D(\eth_udp_inst|crc32_inst|crc_next~5_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [11]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~16_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [11]));
defparam \eth_udp_inst|crc32_inst|crc_data[11] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .coord_z = 3;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .mask = 16'h1122;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[11] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[12] (
	.A(\eth_udp_inst|crc32_inst|crc_next~2_combout ),
	.B(\eth_udp_inst|crc32_inst|crc_data [8]),
	.C(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.D(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [12]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~24_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [12]));
defparam \eth_udp_inst|crc32_inst|crc_data[12] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .coord_y = 8;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .coord_z = 7;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .mask = 16'h0609;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[12] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[13] (
	.A(\eth_udp_inst|crc32_inst|crc_data [9]),
	.B(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.C(\eth_udp_inst|crc32_inst|crc_next~6_combout ),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [13]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~11_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [13]));
defparam \eth_udp_inst|crc32_inst|crc_data[13] .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .coord_z = 6;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[13] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[14] (
	.A(\eth_udp_inst|crc32_inst|crc_data [10]),
	.B(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.C(vcc),
	.D(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [14]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~32_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [14]));
defparam \eth_udp_inst|crc32_inst|crc_data[14] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .coord_y = 8;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .coord_z = 6;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .mask = 16'h1122;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[14] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[15] (
	.A(\eth_udp_inst|crc32_inst|crc_data [11]),
	.B(\eth_udp_inst|crc32_inst|crc_data [31]),
	.C(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [15]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~18_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [15]));
defparam \eth_udp_inst|crc32_inst|crc_data[15] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .coord_z = 1;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .mask = 16'h0609;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[15] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[16] (
	.A(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.B(\eth_udp_inst|crc32_inst|crc_data [12]),
	.C(\eth_udp_inst|crc32_inst|crc_data [28]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [16]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~29_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [16]));
defparam \eth_udp_inst|crc32_inst|crc_data[16] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .coord_y = 8;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .coord_z = 8;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .mask = 16'h1441;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[16] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[17] (
	.A(\eth_udp_inst|crc32_inst|crc_data [13]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.C(\eth_udp_inst|crc32_inst|crc_data [29]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [17]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~15_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [17]));
defparam \eth_udp_inst|crc32_inst|crc_data[17] .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .coord_z = 4;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[17] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[18] (
	.A(\eth_udp_inst|crc32_inst|crc_data [30]),
	.B(\eth_udp_inst|crc32_inst|crc_data [14]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [18]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~35_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [18]));
defparam \eth_udp_inst|crc32_inst|crc_data[18] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .coord_z = 4;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[18] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[19] (
	.A(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.B(\eth_udp_inst|crc32_inst|crc_data [31]),
	.C(\eth_udp_inst|crc32_inst|crc_data [15]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [19]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~21_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [19]));
defparam \eth_udp_inst|crc32_inst|crc_data[19] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .coord_z = 0;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .mask = 16'h1441;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[19] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[1] (
	.A(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.B(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.C(\eth_udp_inst|crc32_inst|crc_data [29]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [1]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~38_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [1]));
defparam \eth_udp_inst|crc32_inst|crc_data[1] .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .coord_z = 15;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .mask = 16'h1441;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[1] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[20] (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|crc32_inst|crc_data [16]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [20]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~26_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [20]));
defparam \eth_udp_inst|crc32_inst|crc_data[20] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .coord_z = 3;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .mask = 16'h00F0;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[20] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[21] (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|crc32_inst|crc_data [17]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [21]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~12_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [21]));
defparam \eth_udp_inst|crc32_inst|crc_data[21] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .coord_z = 15;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .mask = 16'h00F0;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[21] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[22] (
	.A(\eth_udp_inst|crc32_inst|crc_data [28]),
	.B(\eth_udp_inst|crc32_inst|crc_data [18]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [22]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~33_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [22]));
defparam \eth_udp_inst|crc32_inst|crc_data[22] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .coord_z = 0;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[22] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[23] (
	.A(\eth_udp_inst|crc32_inst|crc_data [19]),
	.B(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.C(\eth_udp_inst|crc32_inst|crc_next~6_combout ),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [23]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~19_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [23]));
defparam \eth_udp_inst|crc32_inst|crc_data[23] .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .coord_z = 5;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .mask = 16'h0096;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[23] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[24] (
	.A(\eth_udp_inst|crc32_inst|crc_data [20]),
	.B(\eth_udp_inst|crc32_inst|crc_next~2_combout ),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [24]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~27_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [24]));
defparam \eth_udp_inst|crc32_inst|crc_data[24] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .coord_z = 12;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .mask = 16'h0066;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[24] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[25] (
	.A(\eth_udp_inst|crc32_inst|crc_data [21]),
	.B(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.C(vcc),
	.D(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [25]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~13_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [25]));
defparam \eth_udp_inst|crc32_inst|crc_data[25] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .coord_z = 11;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .mask = 16'h1122;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[25] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[26] (
	.A(\eth_udp_inst|crc32_inst|crc_data [22]),
	.B(\eth_udp_inst|crc32_inst|crc_next~3_combout ),
	.C(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [26]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~34_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [26]));
defparam \eth_udp_inst|crc32_inst|crc_data[26] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .coord_z = 15;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .mask = 16'h0096;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[26] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[27] (
	.A(\eth_udp_inst|crc32_inst|crc_data [23]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.C(\eth_udp_inst|crc32_inst|crc_data [29]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [27]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~20_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [27]));
defparam \eth_udp_inst|crc32_inst|crc_data[27] .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .coord_z = 7;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[27] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[28] (
	.A(\eth_udp_inst|crc32_inst|crc_data [30]),
	.B(\eth_udp_inst|crc32_inst|crc_data [24]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [28]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~37_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [28]));
defparam \eth_udp_inst|crc32_inst|crc_data[28] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .coord_z = 6;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .mask = 16'h0069;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[28] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[29] (
	.A(\eth_udp_inst|crc32_inst|crc_data [25]),
	.B(\eth_udp_inst|crc32_inst|crc_data [31]),
	.C(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [29]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~36_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [29]));
defparam \eth_udp_inst|crc32_inst|crc_data[29] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .coord_z = 6;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .mask = 16'h0609;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[29] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[2] (
	.A(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.C(\eth_udp_inst|crc32_inst|crc_next~2_combout ),
	.D(\eth_udp_inst|crc32_inst|crc_data [28]),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [2]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~40_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [2]));
defparam \eth_udp_inst|crc32_inst|crc_data[2] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .coord_y = 8;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .coord_z = 11;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .mask = 16'h4114;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[2] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[30] (
	.A(\eth_udp_inst|crc32_inst|crc_data [26]),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [30]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~28_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [30]));
defparam \eth_udp_inst|crc32_inst|crc_data[30] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .coord_z = 5;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .mask = 16'h00AA;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[30] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[31] (
	.A(vcc),
	.B(\eth_udp_inst|crc32_inst|crc_data [27]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [31]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~14_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [31]));
defparam \eth_udp_inst|crc32_inst|crc_data[31] .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .coord_z = 10;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .mask = 16'h00CC;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[31] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[3] (
	.A(\eth_udp_inst|crc32_inst|crc_data [29]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.C(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.D(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [3]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~39_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [3]));
defparam \eth_udp_inst|crc32_inst|crc_data[3] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .coord_z = 5;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .mask = 16'h0906;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[3] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[4] (
	.A(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.B(\eth_udp_inst|crc32_inst|crc_data [0]),
	.C(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.D(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [4]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~23_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [4]));
defparam \eth_udp_inst|crc32_inst|crc_data[4] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .coord_y = 8;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .coord_z = 15;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .mask = 16'h1441;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[4] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[5] (
	.A(\eth_udp_inst|crc32_inst|crc_data [1]),
	.B(vcc),
	.C(\eth_udp_inst|crc32_inst|crc_next~5_combout ),
	.D(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [5]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~10_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [5]));
defparam \eth_udp_inst|crc32_inst|crc_data[5] .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .coord_z = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .mask = 16'h005A;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[5] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[6] (
	.A(\eth_udp_inst|crc32_inst|crc_next~2_combout ),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.D(\eth_udp_inst|crc32_inst|crc_data [2]),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [6]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~31_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [6]));
defparam \eth_udp_inst|crc32_inst|crc_data[6] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .coord_y = 8;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .coord_z = 12;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .mask = 16'h050A;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[6] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[7] (
	.A(\eth_udp_inst|crc32_inst|crc_data [3]),
	.B(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.C(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.D(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [7]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~17_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [7]));
defparam \eth_udp_inst|crc32_inst|crc_data[7] .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .coord_z = 13;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .mask = 16'h1221;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[7] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[8] (
	.A(\eth_udp_inst|crc32_inst|crc_data [4]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.D(\eth_udp_inst|crc32_inst|crc_next~5_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [8]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X26_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~22_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [8]));
defparam \eth_udp_inst|crc32_inst|crc_data[8] .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .coord_y = 8;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .coord_z = 2;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .mask = 16'h050A;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[8] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_data[9] (
	.A(vcc),
	.B(\eth_udp_inst|crc32_inst|crc_data [5]),
	.C(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.D(\eth_udp_inst|crc32_inst|crc_next~2_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|crc32_inst|crc_data [9]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|crc32_inst|crc_data[29]~9_combout_X25_Y12_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data~8_combout ),
	.Cout(),
	.Q(\eth_udp_inst|crc32_inst|crc_data [9]));
defparam \eth_udp_inst|crc32_inst|crc_data[9] .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .coord_z = 11;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .mask = 16'h030C;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_data[9] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next[28]~1 (
	.A(\eth_udp_inst|crc32_inst|crc_data [30]),
	.B(\eth_udp_inst|crc32_inst|crc_data [24]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.D(\eth_udp_inst|ip_send_inst|crc_en~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next[28]~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .coord_z = 2;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .mask = 16'h9600;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[28]~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next[29]~0 (
	.A(\eth_udp_inst|crc32_inst|crc_data [25]),
	.B(\eth_udp_inst|ip_send_inst|crc_en~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.D(\eth_udp_inst|crc32_inst|crc_data [31]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next[29]~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .coord_z = 9;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .mask = 16'h8448;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next[29]~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next~2 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.B(\eth_udp_inst|crc32_inst|crc_data [30]),
	.C(\eth_udp_inst|crc32_inst|crc_data [29]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next~2 .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .coord_z = 3;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .mask = 16'h6996;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next~3 (
	.A(vcc),
	.B(\eth_udp_inst|crc32_inst|crc_data [31]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next~3 .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .coord_z = 7;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .mask = 16'h33CC;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next~4 (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|crc32_inst|crc_data [28]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next~4 .coord_x = 22;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .coord_y = 8;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .coord_z = 13;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .mask = 16'h0FF0;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next~5 (
	.A(\eth_udp_inst|crc32_inst|crc_data [29]),
	.B(\eth_udp_inst|crc32_inst|crc_next~3_combout ),
	.C(\eth_udp_inst|crc32_inst|crc_next~4_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next~5_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next~5 .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .coord_z = 12;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .mask = 16'h9669;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~5 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next~6 (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|crc32_inst|crc_data [29]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next~6_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next~6 .coord_x = 21;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .coord_z = 0;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .mask = 16'h0FF0;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~6 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|crc32_inst|crc_next~7 (
	.A(\eth_udp_inst|crc32_inst|crc_data [30]),
	.B(\eth_udp_inst|crc32_inst|crc_data [31]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|crc32_inst|crc_next~7_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|crc32_inst|crc_next~7 .coord_x = 20;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .coord_y = 9;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .coord_z = 8;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .mask = 16'h6996;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .modeMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .ShiftMux = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .BypassEn = 1'b0;
defparam \eth_udp_inst|crc32_inst|crc_next~7 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add13~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt_add [0]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~0 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .mask = 16'h6688;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~10 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~10 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~12 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [6]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~12 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~14 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~14 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~16 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [8]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~16 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~18 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [9]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~18 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~2 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt_add [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~2 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~20 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [10]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~20 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~22 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [11]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~22 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~24 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [12]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~24 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~26 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [13]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~26 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~28 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [14]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~29 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~28 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~28 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~30 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|data_cnt [15]),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~29 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~30_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~30 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .mask = 16'h0FF0;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~30 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add13~4 (
	.A(\eth_udp_inst|ip_send_inst|cnt_add [2]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~4 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~6 (
	.A(\eth_udp_inst|ip_send_inst|cnt_add [3]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~6 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add13~8 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [4]),
	.B(\eth_udp_inst|ip_send_inst|cnt_add [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add13~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add13~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add13~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add13~8 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add13~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .mask = 16'h6688;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~10 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~10 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~12 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~12 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .mask = 16'h964D;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~14 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~14 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~16 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~16 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .mask = 16'h964D;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~18 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~18 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~2 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~2 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~20 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~20 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~22 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~22 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~24 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~24 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .mask = 16'h5AAF;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~26 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~26 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~28 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~28_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~28 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .mask = 16'h0F0F;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~28 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add2~4 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~4 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~6 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~6 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add2~8 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add2~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add2~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add2~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add2~8 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add2~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add3~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add2~24_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add3~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add3~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add3~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .mask = 16'h33CC;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add3~2 (
	.A(\eth_udp_inst|ip_send_inst|Add2~26_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add3~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add3~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add3~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add3~2 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add3~4 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|Add2~28_combout ),
	.Cin(\eth_udp_inst|ip_send_inst|Add3~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add3~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add3~4 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .mask = 16'hF00F;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add3~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add4~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .mask = 16'h6688;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~10 (
	.A(\eth_udp_inst|ip_send_inst|Add2~6_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~10 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~12 (
	.A(\eth_udp_inst|ip_send_inst|Add2~8_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][6]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~12 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~14 (
	.A(\eth_udp_inst|ip_send_inst|Add2~10_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][7]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~14 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~16 (
	.A(\eth_udp_inst|ip_send_inst|Add2~12_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~16 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~18 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][9]~q ),
	.B(\eth_udp_inst|ip_send_inst|Add2~14_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~18 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~2 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][1]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~2 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~20 (
	.A(\eth_udp_inst|ip_send_inst|Add2~16_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][10]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~20 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~22 (
	.A(\eth_udp_inst|ip_send_inst|Add2~18_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][11]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~22 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~24 (
	.A(\eth_udp_inst|ip_send_inst|Add2~20_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][12]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~24 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~26 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][13]~q ),
	.B(\eth_udp_inst|ip_send_inst|Add2~22_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~26 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~28 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][14]~q ),
	.B(\eth_udp_inst|ip_send_inst|Add3~0_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~29 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~28 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~28 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~30 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][15]~q ),
	.B(\eth_udp_inst|ip_send_inst|Add3~2_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~29 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~30_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~31 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~30 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~30 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~32 (
	.A(\eth_udp_inst|ip_send_inst|Add3~4_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~31 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~32_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~33 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~32 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~32 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~34 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~33 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~34_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~34 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .mask = 16'hF0F0;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~34 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add4~4 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][2]~q ),
	.B(\eth_udp_inst|ip_send_inst|Add2~0_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~4 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~6 (
	.A(\eth_udp_inst|ip_send_inst|Add2~2_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][3]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~6 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add4~8 (
	.A(\eth_udp_inst|ip_send_inst|Add2~4_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][4]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add4~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add4~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add4~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add4~8 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add4~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~0_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .mask = 16'h33CC;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~10 (
	.A(\eth_udp_inst|ip_send_inst|Add4~10_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~10 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~12 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~12_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~12 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~14 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~14_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~14 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~16 (
	.A(\eth_udp_inst|ip_send_inst|Add4~16_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~16 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~18 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~18_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~18 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~2 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~2_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~2 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~20 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~20_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~20 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~22 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~22_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~22 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~24 (
	.A(\eth_udp_inst|ip_send_inst|Add4~24_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~24 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~26 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~26_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~26 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~28 (
	.A(\eth_udp_inst|ip_send_inst|Add4~28_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~29 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~28 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .mask = 16'h5AAF;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~28 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~30 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~30_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~29 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~30_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~31 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~30 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~30 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~32 (
	.A(\eth_udp_inst|ip_send_inst|Add4~32_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~31 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~32_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~33 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~32 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~32 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~34 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|Add4~34_combout ),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~33 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~34_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~34 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .mask = 16'h0FF0;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~34 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add5~4 (
	.A(\eth_udp_inst|ip_send_inst|Add4~4_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~4 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~6 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~6_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~6 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add5~8 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add4~8_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add5~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add5~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add5~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add5~8 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .mask = 16'h3CCF;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add5~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~6_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .mask = 16'h33CC;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~10 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~16_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~10 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~12 (
	.A(\eth_udp_inst|ip_send_inst|Add5~18_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~12 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~14 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~20_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~14 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~16 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~22_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~16 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~18 (
	.A(\eth_udp_inst|ip_send_inst|Add5~24_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~18 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~2 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~8_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~2 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~20 (
	.A(\eth_udp_inst|ip_send_inst|Add5~26_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~20 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~22 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~28_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~22 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .mask = 16'hC303;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~24 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~30_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~24 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .mask = 16'h3CCF;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~26 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~32_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~26 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~28 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|Add5~34_combout ),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~28_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~28 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .mask = 16'hF00F;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~28 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add6~4 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~10_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~4 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .mask = 16'h3CCF;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~6 (
	.A(\eth_udp_inst|ip_send_inst|Add5~12_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~6 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add6~8 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~14_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add6~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add6~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add6~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add6~8 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .mask = 16'h3CCF;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add6~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~0 (
	.A(\eth_udp_inst|ip_send_inst|Add5~2_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .mask = 16'h55AA;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~10 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~6_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~10 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~12 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~8_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~12 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~14 (
	.A(\eth_udp_inst|ip_send_inst|Add6~10_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~14 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .mask = 16'hA505;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~16 (
	.A(\eth_udp_inst|ip_send_inst|Add6~12_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~16 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .mask = 16'h5AAF;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~18 (
	.A(\eth_udp_inst|ip_send_inst|Add6~14_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~18 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~2 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~4_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~2 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~20 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~16_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~20 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~22 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~18_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~22 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~24 (
	.A(\eth_udp_inst|ip_send_inst|Add6~20_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~24 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~26 (
	.A(\eth_udp_inst|ip_send_inst|Add6~22_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~26 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~28 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~24_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~29 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~28 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~28 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~30 (
	.A(\eth_udp_inst|ip_send_inst|Add6~26_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~29 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~30_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~31 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~30 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~30 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~32 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|Add6~28_combout ),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~31 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~32_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~32 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .coord_y = 17;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .mask = 16'hF00F;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~32 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add7~4 (
	.A(\eth_udp_inst|ip_send_inst|Add6~0_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~4 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~6 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~2_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~6 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add7~8 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add6~4_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add7~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add7~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add7~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add7~8 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .coord_y = 18;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add7~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~4_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~0 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .mask = 16'h33CC;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~10 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~14_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~10 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~12 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~16_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~12 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~14 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~18_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~14 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~16 (
	.A(\eth_udp_inst|ip_send_inst|Add7~20_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~16 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~18 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~22_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~18 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~2 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~6_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~2 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~20 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~24_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~20 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~22 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~26_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~22 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .mask = 16'hC303;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~24 (
	.A(\eth_udp_inst|ip_send_inst|Add7~28_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~24 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .mask = 16'h5AAF;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~26 (
	.A(\eth_udp_inst|ip_send_inst|Add7~30_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~26 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~28 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~32_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~29 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~28 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~28 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~30 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~29 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~30_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~30 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .mask = 16'hF0F0;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~30 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add8~4 (
	.A(\eth_udp_inst|ip_send_inst|Add7~8_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~4 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .mask = 16'h5AAF;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~6 (
	.A(\eth_udp_inst|ip_send_inst|Add7~10_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~6 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add8~8 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add7~12_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add8~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add8~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add8~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add8~8 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .mask = 16'h3CCF;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add8~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add5~0_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~0_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~1 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .mask = 16'h33CC;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~0 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~10 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~4_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~10_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~11 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~10 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~10 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~12 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~6_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~11 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~12_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~13 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~12 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~12 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~14 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~8_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~15 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~14 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~14 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~16 (
	.A(\eth_udp_inst|ip_send_inst|Add8~10_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~17 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~16 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .mask = 16'h5AAF;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~16 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~18 (
	.A(\eth_udp_inst|ip_send_inst|Add8~12_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~19 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~18 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .mask = 16'hA505;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~18 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~2 (
	.A(\eth_udp_inst|ip_send_inst|Add7~0_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~1 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~2_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~3 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~2 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .mask = 16'hA505;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~2 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~20 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~14_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~21 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~20 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~20 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~22 (
	.A(\eth_udp_inst|ip_send_inst|Add8~16_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~23 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~22 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~22 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~24 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~18_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~23 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~25 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~24 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~24 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~26 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~20_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~25 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~27 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~26 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~26 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~28 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~22_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~27 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~29 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~28 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~28 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~30 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~24_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~29 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~30_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~31 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~30 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~30 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~32 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|Add8~26_combout ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~31 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~32_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~33 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~32 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~32 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~34 (
	.A(\eth_udp_inst|ip_send_inst|Add8~28_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~33 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~34_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~35 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~34 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~34 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~36 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|Add8~30_combout ),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~35 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~36_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~36 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .coord_y = 15;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .mask = 16'hF00F;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~36 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Add9~4 (
	.A(\eth_udp_inst|ip_send_inst|Add7~2_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~4_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~5 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~4 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~4 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~6 (
	.A(\eth_udp_inst|ip_send_inst|Add8~0_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~5 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~6_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~7 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~6 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~6 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Add9~8 (
	.A(\eth_udp_inst|ip_send_inst|Add8~2_combout ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|Add9~7 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Add9~8_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|Add9~9 ),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Add9~8 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .coord_y = 16;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Add9~8 .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|Equal1~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .mask = 16'h1111;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal1~1 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt [4]),
	.C(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal1~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .mask = 16'h0010;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal1~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~0 (
	.A(\eth_udp_inst|ip_send_inst|data_len [10]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|data_cnt [10]),
	.D(\eth_udp_inst|ip_send_inst|data_cnt [9]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .mask = 16'h50A0;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~1 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|data_cnt [3]),
	.D(\eth_udp_inst|ip_send_inst|data_cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .mask = 16'h8000;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~2 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [6]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [4]),
	.C(\eth_udp_inst|ip_send_inst|data_cnt [5]),
	.D(\eth_udp_inst|ip_send_inst|data_cnt [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .mask = 16'h8000;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~3 (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Equal8~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|Equal8~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .mask = 16'hF000;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~4 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [11]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [12]),
	.C(\eth_udp_inst|ip_send_inst|data_cnt [13]),
	.D(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .mask = 16'h0180;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~5 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [14]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [8]),
	.C(\eth_udp_inst|ip_send_inst|data_cnt [15]),
	.D(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~5_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .mask = 16'h0180;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~5 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal8~6 (
	.A(\eth_udp_inst|ip_send_inst|Equal8~3_combout ),
	.B(\eth_udp_inst|ip_send_inst|Equal8~4_combout ),
	.C(\eth_udp_inst|ip_send_inst|Equal8~5_combout ),
	.D(\eth_udp_inst|ip_send_inst|Equal8~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal8~6_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .mask = 16'h8000;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal8~6 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Equal9~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .mask = 16'h0005;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Equal9~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~0 (
	.A(\eth_udp_inst|ip_send_inst|Add13~28_combout ),
	.B(\eth_udp_inst|ip_send_inst|Add13~26_combout ),
	.C(\eth_udp_inst|ip_send_inst|Add13~30_combout ),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .mask = 16'hFEFE;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~1 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|LessThan1~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|Add13~24_combout ),
	.D(\eth_udp_inst|ip_send_inst|Add13~22_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .mask = 16'hFFFC;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~2 (
	.A(\eth_udp_inst|ip_send_inst|Add13~12_combout ),
	.B(\eth_udp_inst|ip_send_inst|data_len [10]),
	.C(\eth_udp_inst|ip_send_inst|Add13~14_combout ),
	.D(\eth_udp_inst|ip_send_inst|Add13~20_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .mask = 16'hB3B2;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~3 (
	.A(\eth_udp_inst|ip_send_inst|Add13~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|data_len [10]),
	.C(\eth_udp_inst|ip_send_inst|Add13~2_combout ),
	.D(\eth_udp_inst|ip_send_inst|Add13~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .mask = 16'hB332;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~4 (
	.A(\eth_udp_inst|ip_send_inst|Add13~6_combout ),
	.B(\eth_udp_inst|ip_send_inst|data_len [10]),
	.C(\eth_udp_inst|ip_send_inst|Add13~8_combout ),
	.D(\eth_udp_inst|ip_send_inst|LessThan1~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .mask = 16'hB020;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~5 (
	.A(\eth_udp_inst|ip_send_inst|LessThan1~4_combout ),
	.B(\eth_udp_inst|ip_send_inst|data_len [10]),
	.C(\eth_udp_inst|ip_send_inst|LessThan1~2_combout ),
	.D(\eth_udp_inst|ip_send_inst|Add13~10_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~5_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .mask = 16'h4CCD;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~5 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~6 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|LessThan1~5_combout ),
	.C(\eth_udp_inst|ip_send_inst|Add13~16_combout ),
	.D(\eth_udp_inst|ip_send_inst|Add13~18_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~6_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .mask = 16'h000C;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~6 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan1~7 (
	.A(\eth_udp_inst|ip_send_inst|LessThan1~6_combout ),
	.B(\eth_udp_inst|ip_send_inst|data_len [10]),
	.C(\eth_udp_inst|ip_send_inst|LessThan1~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|Add13~20_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan1~7_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .mask = 16'h0A0E;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan1~7 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan2~0 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [11]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [12]),
	.C(\eth_udp_inst|ip_send_inst|data_cnt [13]),
	.D(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan2~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .mask = 16'h007F;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan2~1 (
	.A(\eth_udp_inst|ip_send_inst|data_len [10]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [8]),
	.C(\eth_udp_inst|ip_send_inst|Equal8~3_combout ),
	.D(\eth_udp_inst|ip_send_inst|data_cnt [9]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan2~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .mask = 16'h1555;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|LessThan2~2 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [9]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [8]),
	.C(\eth_udp_inst|ip_send_inst|Equal8~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|Equal8~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|LessThan2~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .mask = 16'h0111;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|LessThan2~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux13~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [3]),
	.B(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux13~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .mask = 16'h444C;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux13~1 (
	.A(\eth_udp_inst|ip_send_inst|cnt [3]),
	.B(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux13~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .mask = 16'h0C04;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux13~2 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux13~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .mask = 16'h00CC;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux13~3 (
	.A(\eth_udp_inst|ip_send_inst|cnt [3]),
	.B(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux13~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .mask = 16'h040C;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux13~4 (
	.A(\eth_udp_inst|ip_send_inst|cnt [3]),
	.B(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux13~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .mask = 16'h0C4C;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux13~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux16~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux16~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .mask = 16'h0020;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux16~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux17~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~q ),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux17~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .mask = 16'h44F5;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux17~1 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|Mux17~0_combout ),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux17~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .mask = 16'h8844;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux17~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux20~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux20~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .mask = 16'h50EA;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux20~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux21~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux21~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .mask = 16'h5573;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux21~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux24~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux24~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .mask = 16'hF030;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux24~1 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|Mux24~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux24~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .mask = 16'h320C;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux24~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux25~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux25~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .mask = 16'h0040;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux25~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux27~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux27~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .mask = 16'hFF9D;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux27~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux28~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux28~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .mask = 16'hAFB5;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux28~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux29~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux29~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .mask = 16'h0400;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux29~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux31~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux31~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .mask = 16'hEFBB;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux31~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux32~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[2][11]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux32~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .mask = 16'h1000;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux32~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux33~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.D(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux33~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .mask = 16'hB800;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux33~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux35~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~q ),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux35~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .mask = 16'h5588;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux35~1 (
	.A(\eth_udp_inst|ip_send_inst|cnt [0]),
	.B(\eth_udp_inst|ip_send_inst|Mux35~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux35~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .mask = 16'hE5E4;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux35~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux36~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][15]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux36~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .mask = 16'h5008;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux36~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux37~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][14]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux37~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .mask = 16'hFAF7;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux37~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux39~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][12]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux39~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .mask = 16'h0008;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux39~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux40~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][3]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux40~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .mask = 16'hCA00;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux40~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux41~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][2]~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.D(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux41~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .mask = 16'hB800;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux41~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux43~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][0]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux43~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .mask = 16'hFFB5;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux43~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux44~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][7]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux44~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .mask = 16'h0400;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux44~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux45~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[2][6]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux45~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .mask = 16'h0020;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux45~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|Mux47~0 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.B(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|ip_udp_head[2][4]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|Mux47~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .mask = 16'hC808;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|Mux47~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|always10~0 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always10~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|always10~0 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|always10~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|always10~0 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|always10~0 .mask = 16'h3000;
defparam \eth_udp_inst|ip_send_inst|always10~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always10~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always10~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always10~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always10~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|always3~2 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always3~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|always3~2 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|always3~2 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|always3~2 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|always3~2 .mask = 16'h3000;
defparam \eth_udp_inst|ip_send_inst|always3~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|always3~3 (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt [4]),
	.C(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always3~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|always3~3 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|always3~3 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|always3~3 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|always3~3 .mask = 16'h0030;
defparam \eth_udp_inst|ip_send_inst|always3~3 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|always3~4 (
	.A(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always3~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|always3~4 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|always3~4 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|always3~4 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|always3~4 .mask = 16'h5500;
defparam \eth_udp_inst|ip_send_inst|always3~4 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always3~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|always7~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt [4]),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always7~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|always7~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|always7~0 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|always7~0 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|always7~0 .mask = 16'h0020;
defparam \eth_udp_inst|ip_send_inst|always7~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|always7~1 (
	.A(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.B(\eth_udp_inst|ip_send_inst|always10~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|always7~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always7~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|always7~1 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|always7~1 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|always7~1 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|always7~1 .mask = 16'h0800;
defparam \eth_udp_inst|ip_send_inst|always7~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|always7~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[0] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [16]),
	.B(\eth_udp_inst|ip_send_inst|check_sum [0]),
	.C(\eth_udp_inst|ip_send_inst|Add9~0_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [0]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y15_SIG ),
	.SyncReset(SyncReset_X22_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[0]~17_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[0]~18 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [0]));
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .mask = 16'h6688;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[0] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[10] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [10]),
	.C(\eth_udp_inst|ip_send_inst|Add9~20_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[9]~36 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [10]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y14_SIG ),
	.SyncReset(SyncReset_X22_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[10]~37_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[10]~38 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [10]));
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[10] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[11] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [11]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~22_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[10]~38 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [11]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y14_SIG ),
	.SyncReset(SyncReset_X22_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[11]~39_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[11]~40 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [11]));
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[11] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[12] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [12]),
	.C(\eth_udp_inst|ip_send_inst|Add9~24_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[11]~40 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [12]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y14_SIG ),
	.SyncReset(SyncReset_X22_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[12]~41_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[12]~42 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [12]));
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[12] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[13] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [13]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~26_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[12]~42 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [13]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y14_SIG ),
	.SyncReset(SyncReset_X22_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[13]~43_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[13]~44 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [13]));
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[13] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[14] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [14]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~28_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[13]~44 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [14]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y14_SIG ),
	.SyncReset(SyncReset_X22_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[14]~45_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[14]~46 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [14]));
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[14] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[15] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [15]),
	.C(\eth_udp_inst|ip_send_inst|Add9~30_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[14]~46 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [15]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y14_SIG ),
	.SyncReset(SyncReset_X22_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[15]~48_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[15]~49 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [15]));
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[15] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[16] (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~32_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[15]~49 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [16]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y14_SIG ),
	.SyncReset(SyncReset_X22_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[16]~52_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [16]));
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .mask = 16'h0F0F;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[16] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[17] (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Equal1~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|Add9~34_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [17]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum~51_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [17]));
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .mask = 16'hF000;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[17] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[18] (
	.A(\eth_udp_inst|ip_send_inst|Equal1~1_combout ),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~36_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [18]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum~50_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [18]));
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .mask = 16'hA0A0;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[18] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[1] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [17]),
	.B(\eth_udp_inst|ip_send_inst|check_sum [1]),
	.C(\eth_udp_inst|ip_send_inst|Add9~2_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[0]~18 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [1]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y15_SIG ),
	.SyncReset(SyncReset_X22_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[1]~19_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[1]~20 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [1]));
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .mask = 16'h9617;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[1] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[2] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [18]),
	.B(\eth_udp_inst|ip_send_inst|check_sum [2]),
	.C(\eth_udp_inst|ip_send_inst|Add9~4_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[1]~20 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [2]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y15_SIG ),
	.SyncReset(SyncReset_X22_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[2]~21_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[2]~22 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [2]));
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .mask = 16'h698E;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[2] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[3] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [3]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~6_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[2]~22 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [3]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y15_SIG ),
	.SyncReset(SyncReset_X22_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[3]~23_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[3]~24 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [3]));
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[3] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[4] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [4]),
	.C(\eth_udp_inst|ip_send_inst|Add9~8_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[3]~24 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [4]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y15_SIG ),
	.SyncReset(SyncReset_X22_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[4]~25_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[4]~26 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [4]));
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[4] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[5] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [5]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~10_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[4]~26 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [5]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y15_SIG ),
	.SyncReset(SyncReset_X22_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[5]~27_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[5]~28 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [5]));
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[5] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[6] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [6]),
	.C(\eth_udp_inst|ip_send_inst|Add9~12_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[5]~28 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [6]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y15_SIG ),
	.SyncReset(SyncReset_X22_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[6]~29_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[6]~30 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [6]));
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[6] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[7] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [7]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~14_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[6]~30 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [7]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y15_SIG ),
	.SyncReset(SyncReset_X22_Y15_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y15_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[7]~31_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[7]~32 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [7]));
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[7] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[8] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [8]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~16_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[7]~32 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [8]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y14_SIG ),
	.SyncReset(SyncReset_X22_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[8]~33_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[8]~34 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [8]));
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[8] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[8]~47 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|always3~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[8]~47_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .mask = 16'h1500;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[8]~47 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|check_sum[9] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [9]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|Add9~18_combout ),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|check_sum[8]~34 ),
	.Qin(\eth_udp_inst|ip_send_inst|check_sum [9]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|check_sum[8]~47_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X22_Y14_SIG ),
	.SyncReset(SyncReset_X22_Y14_GND),
	.ShiftData(),
	.SyncLoad(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y14_SIG ),
	.LutOut(\eth_udp_inst|ip_send_inst|check_sum[9]~35_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|check_sum[9]~36 ),
	.Q(\eth_udp_inst|ip_send_inst|check_sum [9]));
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|check_sum[9] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt[0] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[4]~13_combout_X24_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|cnt[4]~11_combout__SyncReset_X24_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X24_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[0]~5_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt[0]~6 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt [0]));
defparam \eth_udp_inst|ip_send_inst|cnt[0] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .mask = 16'h33CC;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[0] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt[1] (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|cnt[0]~6 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[4]~13_combout_X24_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|cnt[4]~11_combout__SyncReset_X24_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X24_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[1]~7_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt[1]~8 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt [1]));
defparam \eth_udp_inst|ip_send_inst|cnt[1] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[1] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt[2] (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|cnt[1]~8 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt [2]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[4]~13_combout_X24_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|cnt[4]~11_combout__SyncReset_X24_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X24_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[2]~9_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt[2]~10 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt [2]));
defparam \eth_udp_inst|ip_send_inst|cnt[2] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[2] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt[3] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|cnt[2]~10 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt [3]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[4]~13_combout_X24_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|cnt[4]~11_combout__SyncReset_X24_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X24_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[3]~14_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt[3]~15 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt [3]));
defparam \eth_udp_inst|ip_send_inst|cnt[3] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[3] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt[4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt [4]),
	.Cin(\eth_udp_inst|ip_send_inst|cnt[3]~15 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt [4]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt[4]~13_combout_X24_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|cnt[4]~11_combout__SyncReset_X24_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X24_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[4]~16_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|cnt [4]));
defparam \eth_udp_inst|ip_send_inst|cnt[4] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .mask = 16'hF00F;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt[4] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt[4]~11 (
	.A(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.B(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.C(\eth_udp_inst|ip_send_inst|always3~2_combout ),
	.D(\eth_udp_inst|ip_send_inst|always3~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[4]~11_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|cnt[4]~11 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~11 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~11 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~11 .mask = 16'hF222;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~11 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~11 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~11 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~11 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~11 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt[4]~12 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[4]~12_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|cnt[4]~12 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~12 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~12 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~12 .mask = 16'h7FFF;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~12 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~12 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt[4]~13 (
	.A(\eth_udp_inst|ip_send_inst|cnt[4]~12_combout ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.D(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt[4]~13_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|cnt[4]~13 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~13 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~13 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~13 .mask = 16'hF4F7;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~13 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~13 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~13 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~13 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt[4]~13 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_add[0] (
	.A(\eth_udp_inst|ip_send_inst|cnt_add [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_add [0]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X26_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[0]~5_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt_add[0]~6 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt_add [0]));
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .mask = 16'h55AA;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[0] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt_add[1] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt_add [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|cnt_add[0]~6 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_add [1]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X26_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[1]~7_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt_add[1]~8 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt_add [1]));
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[1] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt_add[2] (
	.A(\eth_udp_inst|ip_send_inst|cnt_add [2]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|cnt_add[1]~8 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_add [2]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X26_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[2]~9_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt_add[2]~10 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt_add [2]));
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[2] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt_add[3] (
	.A(\eth_udp_inst|ip_send_inst|cnt_add [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|cnt_add[2]~10 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_add [3]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X26_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[3]~11_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|cnt_add[3]~12 ),
	.Q(\eth_udp_inst|ip_send_inst|cnt_add [3]));
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[3] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|cnt_add[4] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt_add [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|cnt_add[3]~12 ),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_add [4]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout_X26_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y16_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y16_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y16_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[4]~13_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|cnt_add [4]));
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .mask = 16'hC3C3;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_add[4]~15 (
	.A(\eth_udp_inst|ip_send_inst|Equal8~6_combout ),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[4]~15_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .mask = 16'h0A0A;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_add[4]~15 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_send_bit[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout_X25_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_send_bit~5_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]));
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .mask = 16'h0F00;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[0] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_send_bit[1] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout_X25_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_send_bit~4_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]));
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .mask = 16'h3C00;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[1] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_send_bit[2] (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1_combout ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout_X25_Y13_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y13_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_send_bit~2_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]));
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .mask = 16'h28A0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 (
	.A(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.B(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .mask = 16'h1111;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.C(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .mask = 16'h72FA;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|cnt_send_bit[2]~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|crc_clr (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|send_end~q ),
	.D(\eth_udp_inst|ip_send_inst|crc_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|crc_clr~q ),
	.Clk(\clk_25m~clkctrl_outclk_X25_Y12_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y12_SIG ),
	.SyncReset(SyncReset_X25_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y12_VCC),
	.LutOut(\eth_udp_inst|crc32_inst|crc_data[29]~9_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|crc_clr~q ));
defparam \eth_udp_inst|ip_send_inst|crc_clr .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|crc_clr .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|crc_clr .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|crc_clr .mask = 16'hFFF0;
defparam \eth_udp_inst|ip_send_inst|crc_clr .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|crc_clr .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|crc_clr .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|crc_clr .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|crc_clr .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|crc_en (
	.A(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|crc_en~q ),
	.Clk(\clk_25m~clkctrl_outclk_X25_Y15_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always13~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|crc_en~q ));
defparam \eth_udp_inst|ip_send_inst|crc_en .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|crc_en .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|crc_en .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|crc_en .mask = 16'hFFFA;
defparam \eth_udp_inst|ip_send_inst|crc_en .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|crc_en .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|crc_en .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|crc_en .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|crc_en .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[0] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [0]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[0]~16_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[0]~17 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [0]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .mask = 16'h55AA;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[0] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[10] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [10]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[9]~35 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [10]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[10]~36_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[10]~37 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [10]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[10]~41 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.C(\eth_udp_inst|ip_send_inst|data_cnt[9]~40_combout ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .mask = 16'hC040;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[10]~41 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[11] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [11]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[10]~37 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [11]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[11]~42_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[11]~43 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [11]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[11] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[12] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [12]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[11]~43 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [12]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[12]~44_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[12]~45 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [12]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[12] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[13] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [13]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[12]~45 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [13]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[13]~46_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[13]~47 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [13]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[13] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[14] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [14]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[13]~47 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [14]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[14]~48_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[14]~49 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [14]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[14] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[15] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [15]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[14]~49 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [15]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[15]~50_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [15]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .mask = 16'h5A5A;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[15] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[1] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[0]~17 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [1]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[1]~18_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[1]~19 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [1]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[1] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[2] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[1]~19 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [2]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[2]~20_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[2]~21 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [2]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[2] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[3] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[2]~21 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [3]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[3]~22_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[3]~23 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [3]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[3] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[4] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[3]~23 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [4]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[4]~24_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[4]~25 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [4]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[4] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[5] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [5]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[4]~25 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [5]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[5]~26_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[5]~27 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [5]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[5] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[6] (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[5]~27 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [6]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[6]~28_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[6]~29 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [6]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[6] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[7] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[6]~29 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [7]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[7]~30_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[7]~31 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [7]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[7] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[8] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [8]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[7]~31 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [8]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[8]~32_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[8]~33 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [8]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[8] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[9] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|data_cnt [9]),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|data_cnt[8]~33 ),
	.Qin(\eth_udp_inst|ip_send_inst|data_cnt [9]),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|data_cnt[10]~41_combout_X26_Y15_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y15_SIG ),
	.SyncReset(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X26_Y15_GND),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[9]~34_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|data_cnt[9]~35 ),
	.Q(\eth_udp_inst|ip_send_inst|data_cnt [9]));
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[9]~38 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [10]),
	.B(\eth_udp_inst|ip_send_inst|LessThan2~2_combout ),
	.C(\eth_udp_inst|ip_send_inst|Equal8~4_combout ),
	.D(\eth_udp_inst|ip_send_inst|LessThan2~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[9]~38_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~38 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~38 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~38 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~38 .mask = 16'hF0D0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~38 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~38 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~38 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~38 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~38 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[9]~39 (
	.A(\eth_udp_inst|ip_send_inst|data_cnt [15]),
	.B(\eth_udp_inst|ip_send_inst|data_cnt[9]~38_combout ),
	.C(\eth_udp_inst|ip_send_inst|LessThan2~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[9]~39_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~39 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~39 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~39 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~39 .mask = 16'h5402;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~39 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~39 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~39 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~39 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~39 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|data_cnt[9]~40 (
	.A(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.B(\eth_udp_inst|ip_send_inst|data_cnt[9]~39_combout ),
	.C(\eth_udp_inst|ip_send_inst|data_cnt [14]),
	.D(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|data_cnt[9]~40_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~40 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~40 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~40 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~40 .mask = 16'hAEBF;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~40 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~40 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~40 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~40 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_cnt[9]~40 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|data_len[10] (
	.A(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.B(\eth_udp_inst|ip_send_inst|send_en_r~q ),
	.C(vcc),
	.D(\LessThan0~0_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|data_len [10]),
	.Clk(\clk_25m~clkctrl_outclk_X24_Y16_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|data_len[10]~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|data_len [10]));
defparam \eth_udp_inst|ip_send_inst|data_len[10] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .mask = 16'hF1F0;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|data_len[10] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data[0] (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~23_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~35_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~42_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.Clk(\clk_25m~clkctrl_outclk_X23_Y16_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~43_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|eth_tx_data [0]));
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .mask = 16'hFEAA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[0] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data[1] (
	.A(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.B(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~90_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~68_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.Clk(\clk_25m~clkctrl_outclk_X23_Y16_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~91_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|eth_tx_data [1]));
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .mask = 16'h3210;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[1] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data[2] (
	.A(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.B(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~19_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.Clk(\clk_25m~clkctrl_outclk_X23_Y16_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~20_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|eth_tx_data [2]));
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .mask = 16'hFF88;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[2] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data[3] (
	.A(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~65_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~64_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.Clk(\clk_25m~clkctrl_outclk_X23_Y16_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~66_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|eth_tx_data [3]));
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .mask = 16'hF4F0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data[3] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~0 (
	.A(\eth_udp_inst|ip_send_inst|Mux13~2_combout ),
	.B(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|Mux13~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .mask = 16'hF2C2;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~1 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|Mux13~3_combout ),
	.C(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|Mux13~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~1_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .mask = 16'hDA8A;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~1 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~10 (
	.A(\eth_udp_inst|crc32_inst|crc_data [21]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~9_combout ),
	.C(\eth_udp_inst|crc32_inst|crc_data [17]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~10_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .mask = 16'hE2CC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~10 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~11 (
	.A(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~8_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~10_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~11_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .mask = 16'h88A0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~11 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~12 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~11_combout ),
	.C(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.D(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~12_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .mask = 16'h00CE;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~12 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~13 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\cmos1_fifo_inst|q [26]),
	.D(\cmos1_fifo_inst|q [18]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~13_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .mask = 16'hB9A8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~13 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~14 (
	.A(\cmos1_fifo_inst|q [30]),
	.B(\cmos1_fifo_inst|q [22]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~13_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~14_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .mask = 16'hACF0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~14 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~15 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(\cmos1_fifo_inst|q [2]),
	.C(\cmos1_fifo_inst|q [6]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~15_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .mask = 16'hAAE4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~15 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~16 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~15_combout ),
	.B(\cmos1_fifo_inst|q [14]),
	.C(\cmos1_fifo_inst|q [10]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~16_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .mask = 16'hD8AA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~16 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~17 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~16_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~14_combout ),
	.D(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~17_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .mask = 16'hE400;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~17 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~18 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~17_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~6_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~12_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~18_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .mask = 16'hF3F2;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~18 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~19 (
	.A(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.B(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~18_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~19_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .mask = 16'h3120;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~19 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~2 (
	.A(\eth_udp_inst|ip_send_inst|Mux33~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.C(\eth_udp_inst|ip_send_inst|Mux41~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .mask = 16'hCCE2;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~21 (
	.A(\eth_udp_inst|ip_send_inst|cnt [3]),
	.B(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~21_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .mask = 16'hF2B0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~21 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~22 (
	.A(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|cnt [3]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~21_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~22_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .mask = 16'h022A;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~22 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~23 (
	.A(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.B(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~22_combout ),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~23_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .mask = 16'hA8A8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~23 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~24 (
	.A(\cmos1_fifo_inst|q [16]),
	.B(\cmos1_fifo_inst|q [20]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~24_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .mask = 16'hFC0A;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~24 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~25 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\cmos1_fifo_inst|q [28]),
	.C(\cmos1_fifo_inst|q [24]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~24_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~25_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .mask = 16'hDDA0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~25 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~26 (
	.A(\cmos1_fifo_inst|q [0]),
	.B(\cmos1_fifo_inst|q [4]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~26_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .mask = 16'hFC0A;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~26 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~27 (
	.A(\cmos1_fifo_inst|q [8]),
	.B(\cmos1_fifo_inst|q [12]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~26_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~27_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .mask = 16'hCFA0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~27 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~28 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.B(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~27_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~25_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~28_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .mask = 16'hC840;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~28 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~29 (
	.A(\eth_udp_inst|crc32_inst|crc_data [7]),
	.B(\eth_udp_inst|crc32_inst|crc_data [15]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~29_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .mask = 16'hF0AC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~29 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~3 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(\eth_udp_inst|ip_send_inst|Mux45~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|Mux37~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .mask = 16'hDD0A;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~30 (
	.A(\eth_udp_inst|crc32_inst|crc_data [3]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~29_combout ),
	.C(\eth_udp_inst|crc32_inst|crc_data [11]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~30_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .mask = 16'hB8CC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~30 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~31 (
	.A(\eth_udp_inst|ip_send_inst|crc_en~q ),
	.B(\eth_udp_inst|crc32_inst|crc_data [27]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~31_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .mask = 16'hFC0D;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~31 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~32 (
	.A(\eth_udp_inst|crc32_inst|crc_data [23]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~31_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|crc32_inst|crc_data [19]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~32_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .mask = 16'hEC2C;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~32 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~33 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.B(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~32_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~30_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~33_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .mask = 16'hC840;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~33 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~34 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.B(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.C(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~33_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~34_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .mask = 16'h3302;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~34 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~35 (
	.A(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~34_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~28_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~35_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .mask = 16'h5550;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~35 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~36 (
	.A(\eth_udp_inst|ip_send_inst|Mux35~1_combout ),
	.B(\eth_udp_inst|ip_send_inst|Mux39~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~36_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .mask = 16'hFC0A;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~36 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~37 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~36_combout ),
	.B(\eth_udp_inst|ip_send_inst|Mux47~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|Mux43~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~37_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .mask = 16'h8ADA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~37 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~38 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~38_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .mask = 16'hDFAA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~38 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~39 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~q ),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~39_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .mask = 16'h8D00;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~39 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~4 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(\eth_udp_inst|ip_send_inst|Mux17~1_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|Mux21~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .mask = 16'hAEA4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~40 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~38_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~39_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~40_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .mask = 16'h8A89;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~40 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~41 (
	.A(\eth_udp_inst|ip_send_inst|Mux27~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~40_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|Mux31~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~41_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .mask = 16'h1CDC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~41 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~42 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~37_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~41_combout ),
	.C(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~42_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .mask = 16'hA0C0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~42 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~44 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~44_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .mask = 16'h00D5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~44 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~45 (
	.A(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|cnt [2]),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~45_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .mask = 16'h1038;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~45 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~46 (
	.A(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~44_combout ),
	.C(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~45_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~46_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .mask = 16'hA080;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~46 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~47 (
	.A(\eth_udp_inst|ip_send_inst|Mux40~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.D(\eth_udp_inst|ip_send_inst|Mux32~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~47_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .mask = 16'hCBC8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~47 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~48 (
	.A(\eth_udp_inst|ip_send_inst|Mux44~0_combout ),
	.B(\eth_udp_inst|ip_send_inst|Mux36~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~47_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~48_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .mask = 16'hAFC0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~48 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~49 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.C(\eth_udp_inst|ip_send_inst|Mux20~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|Mux16~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~49_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .mask = 16'hB9A8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~49 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~5 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~4_combout ),
	.C(\eth_udp_inst|ip_send_inst|Mux29~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|Mux25~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~5_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .mask = 16'hE6C4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~5 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~50 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~49_combout ),
	.B(\eth_udp_inst|ip_send_inst|Mux24~1_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|Mux28~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~50_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .mask = 16'h4AEA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~50 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~51 (
	.A(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~50_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~48_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~51_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .mask = 16'hA820;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~51 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~52 (
	.A(\eth_udp_inst|crc32_inst|crc_data [4]),
	.B(\eth_udp_inst|crc32_inst|crc_data [12]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~52_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .coord_y = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .mask = 16'hF0AC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~52 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~53 (
	.A(\eth_udp_inst|crc32_inst|crc_data [8]),
	.B(\eth_udp_inst|crc32_inst|crc_data [0]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~52_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~53_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .coord_y = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .mask = 16'hCAF0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~53 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~54 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(\eth_udp_inst|crc32_inst|crc_data [24]),
	.C(\eth_udp_inst|crc32_inst|crc_next[28]~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~54_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .mask = 16'hAA8D;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~54 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~55 (
	.A(\eth_udp_inst|crc32_inst|crc_data [16]),
	.B(\eth_udp_inst|crc32_inst|crc_data [20]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~54_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~55_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .mask = 16'hACF0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~55 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~56 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~55_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~53_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~56_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .mask = 16'hC088;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~56 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~57 (
	.A(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.C(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~56_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~57_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .mask = 16'h5504;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~57 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~58 (
	.A(\cmos1_fifo_inst|q [27]),
	.B(\cmos1_fifo_inst|q [19]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~58_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .mask = 16'hF0AC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~58 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~59 (
	.A(\cmos1_fifo_inst|q [31]),
	.B(\cmos1_fifo_inst|q [23]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~58_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~59_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .mask = 16'hACF0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~59 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~6 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~3_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~5_combout ),
	.C(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~6_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .mask = 16'hA0C0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~6 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~60 (
	.A(\cmos1_fifo_inst|q [3]),
	.B(\cmos1_fifo_inst|q [7]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~60_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .mask = 16'hFC0A;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~60 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~61 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~60_combout ),
	.B(\cmos1_fifo_inst|q [11]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\cmos1_fifo_inst|q [15]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~61_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .mask = 16'hEA4A;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~61 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~62 (
	.A(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~61_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~59_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~62_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .mask = 16'hA820;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~62 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~63 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~62_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~51_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~57_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~63_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .mask = 16'hF3F2;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~63 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~65 (
	.A(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.B(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~65_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .mask = 16'h8000;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~65 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~67 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|Mux13~3_combout ),
	.C(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|Mux13~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~67_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .mask = 16'hADA8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~67 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~68 (
	.A(\eth_udp_inst|ip_send_inst|Mux13~2_combout ),
	.B(\eth_udp_inst|ip_send_inst|Mux13~4_combout ),
	.C(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~67_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~68_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .mask = 16'hCFA0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~68 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~69 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[2][13]~q ),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[2][5]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~69_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .mask = 16'hE4AA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~69 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~7 (
	.A(\eth_udp_inst|crc32_inst|crc_data [13]),
	.B(\eth_udp_inst|crc32_inst|crc_data [5]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~7_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .mask = 16'hF0CA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~7 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~70 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[2][1]~q ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~69_combout ),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[2][9]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~70_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .mask = 16'hCCB8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~70 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~71 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~70_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~71_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .mask = 16'h5DF8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~71 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~72 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~71_combout ),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|cnt [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~72_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .mask = 16'h05A0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~72 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~73 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~73_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .mask = 16'hACAC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~73 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~74 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~74_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .mask = 16'hBA00;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~74 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~75 (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~75_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .mask = 16'h3DCC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~75 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~76 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~75_combout ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~q ),
	.C(\eth_udp_inst|ip_send_inst|cnt [0]),
	.D(\eth_udp_inst|ip_send_inst|cnt [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~76_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .mask = 16'h0AD0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~76 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~77 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~75_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~74_combout ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~76_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~73_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~77_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .mask = 16'hD0C0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~77 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~78 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~77_combout ),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~72_combout ),
	.C(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~78_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .mask = 16'hC0A0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~78 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~79 (
	.A(\cmos1_fifo_inst|q [25]),
	.B(\cmos1_fifo_inst|q [17]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~79_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .mask = 16'hF0AC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~79 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~8 (
	.A(\eth_udp_inst|crc32_inst|crc_data [1]),
	.B(\eth_udp_inst|crc32_inst|crc_data [9]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~7_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~8_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .mask = 16'hACF0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~8 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~80 (
	.A(\cmos1_fifo_inst|q [21]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~79_combout ),
	.C(\cmos1_fifo_inst|q [29]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~80_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .mask = 16'hE2CC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~80 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~81 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\cmos1_fifo_inst|q [5]),
	.D(\cmos1_fifo_inst|q [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~81_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .mask = 16'hD9C8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~81 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~82 (
	.A(\cmos1_fifo_inst|q [9]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~81_combout ),
	.C(\cmos1_fifo_inst|q [13]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~82_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .mask = 16'hE2CC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~82 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~83 (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.B(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~82_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~80_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~83_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .mask = 16'hC840;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~83 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~84 (
	.A(\eth_udp_inst|crc32_inst|crc_data [14]),
	.B(\eth_udp_inst|crc32_inst|crc_data [6]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~84_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .coord_y = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .mask = 16'hF0CA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~84 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~85 (
	.A(\eth_udp_inst|crc32_inst|crc_data [10]),
	.B(\eth_udp_inst|ip_send_inst|eth_tx_data~84_combout ),
	.C(\eth_udp_inst|crc32_inst|crc_data [2]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~85_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .coord_y = 8;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .mask = 16'hE2CC;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~85 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~86 (
	.A(\eth_udp_inst|crc32_inst|crc_data [26]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.D(\eth_udp_inst|ip_send_inst|crc_en~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~86_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .mask = 16'hE2E3;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~86 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~87 (
	.A(\eth_udp_inst|crc32_inst|crc_data [22]),
	.B(\eth_udp_inst|crc32_inst|crc_data [18]),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~86_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~87_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .coord_x = 22;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .mask = 16'hCAF0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~87 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~88 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~87_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~85_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~88_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .mask = 16'hC088;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~88 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~89 (
	.A(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.B(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~88_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~89_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .mask = 16'h5150;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~89 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~9 (
	.A(\eth_udp_inst|crc32_inst|crc_data [25]),
	.B(\eth_udp_inst|crc32_inst|crc_next[29]~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~9_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .coord_y = 9;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .mask = 16'hFA03;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~9 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_data~90 (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~78_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data~83_combout ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~89_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~90_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .coord_y = 11;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .mask = 16'hBBBA;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_data~90 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|eth_tx_en (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|eth_tx_en~q ),
	.Clk(\clk_25m~clkctrl_outclk_X25_Y15_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always11~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|eth_tx_en~q ));
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .mask = 16'h00F0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|eth_tx_en .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] (
	.A(\eth_udp_inst|ip_send_inst|data_len [10]),
	.B(\eth_udp_inst|ip_send_inst|always3~4_combout ),
	.C(vcc),
	.D(\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ),
	.Clk(\clk_25m~clkctrl_outclk_X25_Y15_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~18_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[0][10]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .mask = 16'hF0B8;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[0][10] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] (
	.A(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~q ),
	.Clk(\clk_25m~clkctrl_outclk_X25_Y15_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~53_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .mask = 16'hA5F0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][16] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~q ),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][16]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~21_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~22 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .mask = 16'h6688;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][17] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][17]~22 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~23_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~24 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][18] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][18]~24 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~25_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~26 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][19] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][19]~26 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~27_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~28 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][20] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][20]~28 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~29_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~30 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][21] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][21]~30 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~31_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~32 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .coord_z = 6;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .mask = 16'h5A5F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][22] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][22]~32 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~33_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~34 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][23] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][23]~34 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~35_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~36 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .coord_z = 8;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][24] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][24]~36 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~37_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~38 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .mask = 16'hC30C;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][25] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][25]~38 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~39_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~40 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][26] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][26]~40 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~41_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~42 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][27] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][27]~42 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~43_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~44 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][28] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][28]~44 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~45_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~46 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .mask = 16'hA50A;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][29] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][29]~46 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~47_combout ),
	.Cout(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~48 ),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .mask = 16'h3C3F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][30] .CarryEnb = 1'b0;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] (
	.A(\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][30]~48 ),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|always3~4_combout_X21_Y14_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X21_Y14_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~58_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[1][31]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .mask = 16'hA5A5;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .modeMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[1][31] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] (
	.A(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.B(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.C(\eth_udp_inst|ip_send_inst|check_sum [0]),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][0]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X25_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X25_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~49_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][0]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .mask = 16'h0D0D;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][0] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [10]),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][10]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~19_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][10]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .mask = 16'h3033;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][10] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [11]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][11]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~56_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][11]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .mask = 16'h5055;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][11] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [12]),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][12]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~50_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][12]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .mask = 16'h3033;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][12] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [13]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][13]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~62_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][13]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .mask = 16'h5055;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][13] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [14]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][14]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~15_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][14]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .mask = 16'h5055;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][14] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.C(\eth_udp_inst|ip_send_inst|check_sum [15]),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][15]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X25_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X25_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~54_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][15]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .mask = 16'h0C0F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][15] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [1]),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][1]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~60_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][1]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .mask = 16'h3033;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][1] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [2]),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][2]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~17_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][2]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .coord_z = 0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .mask = 16'h3033;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][2] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [3]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][3]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~55_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][3]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .coord_z = 2;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .mask = 16'h5055;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][3] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.C(\eth_udp_inst|ip_send_inst|check_sum [4]),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][4]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X25_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X25_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~52_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][4]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .mask = 16'h0C0F;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][4] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [5]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][5]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~63_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][5]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .coord_z = 5;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .mask = 16'h5055;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][5] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] (
	.A(vcc),
	.B(\eth_udp_inst|ip_send_inst|check_sum [6]),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][6]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~20_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][6]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .coord_z = 1;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .mask = 16'h3033;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][6] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [7]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][7]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y15_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y15_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~57_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][7]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .mask = 16'h5055;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][7] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [8]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~51_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .mask = 16'h5055;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 (
	.A(\eth_udp_inst|ip_send_inst|always3~2_combout ),
	.B(\eth_udp_inst|ip_send_inst|always3~4_combout ),
	.C(\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.D(\eth_udp_inst|ip_send_inst|always3~3_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .mask = 16'h0E0C;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] (
	.A(\eth_udp_inst|ip_send_inst|check_sum [9]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|ip_udp_head[2][9]~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|ip_udp_head[2][8]~16_combout_X22_Y14_SIG_SIG ),
	.AsyncReset(AsyncReset_X22_Y14_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|ip_udp_head~61_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|ip_udp_head[2][9]~q ));
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .coord_y = 13;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .mask = 16'h5055;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|ip_udp_head[2][9] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|packet_head[7][7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ),
	.Clk(\clk_25m~clkctrl_outclk_X23_Y16_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|packet_head[7][7]~feeder_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|packet_head[7][7]~q ));
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .mask = 16'hFFFF;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|packet_head[7][7] .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|read_data_req (
	.A(\eth_udp_inst|ip_send_inst|always7~1_combout ),
	.B(\eth_udp_inst|ip_send_inst|always10~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|Equal8~6_combout ),
	.D(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|read_data_req~q ),
	.Clk(\clk_25m~clkctrl_outclk_X25_Y15_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X25_Y15_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|read_data_req~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|read_data_req~q ));
defparam \eth_udp_inst|ip_send_inst|read_data_req .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|read_data_req .coord_y = 14;
defparam \eth_udp_inst|ip_send_inst|read_data_req .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|read_data_req .mask = 16'hAEAA;
defparam \eth_udp_inst|ip_send_inst|read_data_req .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|read_data_req .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|read_data_req .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|read_data_req .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|read_data_req .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|send_en_r (
	.A(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~14_combout ),
	.B(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~18_combout ),
	.C(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~16_combout ),
	.D(\cmos1_fifo_inst|dcfifo_mixed_widths_component|auto_generated|op_1~12_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|send_en_r~q ),
	.Clk(\clk_25m~clkctrl_outclk_X24_Y16_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\LessThan0~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|send_en_r~q ));
defparam \eth_udp_inst|ip_send_inst|send_en_r .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|send_en_r .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|send_en_r .coord_z = 10;
defparam \eth_udp_inst|ip_send_inst|send_en_r .mask = 16'hFCEC;
defparam \eth_udp_inst|ip_send_inst|send_en_r .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_en_r .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_en_r .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_en_r .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_en_r .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|send_end (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.C(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|send_end~q ),
	.Clk(\clk_25m~clkctrl_outclk_X24_Y12_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|always16~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|send_end~q ));
defparam \eth_udp_inst|ip_send_inst|send_end .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|send_end .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|send_end .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|send_end .mask = 16'h8000;
defparam \eth_udp_inst|ip_send_inst|send_end .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_end .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_end .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_end .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|send_end .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.CHECK_SUM (
	.A(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X26_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ));
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .mask = 16'h5555;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.CHECK_SUM .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.CRC (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [2]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit [1]),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X24_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ),
	.SyncReset(SyncReset_X24_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X24_Y16_VCC),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~5_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.CRC~q ));
defparam \eth_udp_inst|ip_send_inst|state.CRC .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|state.CRC .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|state.CRC .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|state.CRC .mask = 16'hA000;
defparam \eth_udp_inst|ip_send_inst|state.CRC .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.CRC .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.CRC .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.CRC .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.CRC .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.ETH_HEAD (
	.A(\eth_udp_inst|ip_send_inst|eth_tx_data~46_combout ),
	.B(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.C(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data~63_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(SyncReset_X23_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y16_VCC),
	.LutOut(\eth_udp_inst|ip_send_inst|eth_tx_data~64_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ));
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .coord_z = 11;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .mask = 16'h2322;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.ETH_HEAD .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.IDLE (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.D(vcc),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X26_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X26_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|state.IDLE~0_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.IDLE~q ));
defparam \eth_udp_inst|ip_send_inst|state.IDLE .coord_x = 19;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .coord_z = 13;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .mask = 16'h0F0F;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.IDLE .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD (
	.A(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.B(\eth_udp_inst|ip_send_inst|state.CRC~q ),
	.C(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~0_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(SyncReset_X23_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y16_VCC),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_send_bit[2]~3_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ));
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .coord_z = 15;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .mask = 16'hFEFF;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.PACKET_HEAD (
	.A(\eth_udp_inst|ip_send_inst|cnt [3]),
	.B(\eth_udp_inst|ip_send_inst|cnt [1]),
	.C(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.D(\eth_udp_inst|ip_send_inst|state.ETH_HEAD~q ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X23_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X23_Y16_SIG ),
	.SyncReset(SyncReset_X23_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X23_Y16_VCC),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~1_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.PACKET_HEAD~q ));
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .mask = 16'h6240;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.PACKET_HEAD .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|state.SEND_DATA (
	.A(\eth_udp_inst|ip_send_inst|cnt_add[4]~15_combout ),
	.B(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.C(\eth_udp_inst|ip_send_inst|state.IP_UDP_HEAD~q ),
	.D(\eth_udp_inst|ip_send_inst|LessThan1~7_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.Clk(\clk_25m~clkctrl_outclk__eth_udp_inst|ip_send_inst|sw_en~q_X24_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ),
	.SyncReset(SyncReset_X24_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X24_Y16_VCC),
	.LutOut(\eth_udp_inst|ip_send_inst|cnt_add[4]~16_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ));
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .coord_z = 7;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .mask = 16'hE0C0;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .FeedbackMux = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .BypassEn = 1'b1;
defparam \eth_udp_inst|ip_send_inst|state.SEND_DATA .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|sw_en (
	.A(\eth_udp_inst|ip_send_inst|cnt_send_bit [0]),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|sw_en~6_combout ),
	.D(\eth_udp_inst|ip_send_inst|sw_en~4_combout ),
	.Cin(),
	.Qin(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Clk(\clk_25m~clkctrl_outclk_X24_Y16_SIG_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X24_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~7_combout ),
	.Cout(),
	.Q(\eth_udp_inst|ip_send_inst|sw_en~q ));
defparam \eth_udp_inst|ip_send_inst|sw_en .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|sw_en .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|sw_en .coord_z = 4;
defparam \eth_udp_inst|ip_send_inst|sw_en .mask = 16'hFF50;
defparam \eth_udp_inst|ip_send_inst|sw_en .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|sw_en~0 (
	.A(\eth_udp_inst|ip_send_inst|cnt [1]),
	.B(\eth_udp_inst|ip_send_inst|state.CHECK_SUM~q ),
	.C(\eth_udp_inst|ip_send_inst|Equal1~0_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~0_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .mask = 16'h0080;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~0 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|sw_en~2 (
	.A(\eth_udp_inst|ip_send_inst|cnt [2]),
	.B(\eth_udp_inst|ip_send_inst|cnt [0]),
	.C(\eth_udp_inst|ip_send_inst|sw_en~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|Equal9~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~2_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .coord_z = 3;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .mask = 16'h8000;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~2 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|sw_en~3 (
	.A(\eth_udp_inst|ip_send_inst|sw_en~2_combout ),
	.B(\eth_udp_inst|ip_send_inst|sw_en~0_combout ),
	.C(\eth_udp_inst|ip_send_inst|always7~1_combout ),
	.D(\eth_udp_inst|ip_send_inst|cnt [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~3_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .coord_x = 21;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .coord_y = 10;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .coord_z = 9;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .mask = 16'hF0FE;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~3 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|sw_en~4 (
	.A(\eth_udp_inst|ip_send_inst|state.IDLE~q ),
	.B(\eth_udp_inst|ip_send_inst|send_en_r~q ),
	.C(\eth_udp_inst|ip_send_inst|sw_en~3_combout ),
	.D(\LessThan0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~4_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .coord_z = 14;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .mask = 16'hF1F0;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~4 .CarryEnb = 1'b1;

alta_slice \eth_udp_inst|ip_send_inst|sw_en~6 (
	.A(\eth_udp_inst|ip_send_inst|state.SEND_DATA~q ),
	.B(\eth_udp_inst|ip_send_inst|Equal8~6_combout ),
	.C(\eth_udp_inst|ip_send_inst|sw_en~5_combout ),
	.D(\eth_udp_inst|ip_send_inst|LessThan1~7_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\eth_udp_inst|ip_send_inst|sw_en~6_combout ),
	.Cout(),
	.Q());
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .coord_x = 20;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .coord_y = 12;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .coord_z = 12;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .mask = 16'hF0F8;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .modeMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .FeedbackMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .ShiftMux = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .BypassEn = 1'b0;
defparam \eth_udp_inst|ip_send_inst|sw_en~6 .CarryEnb = 1'b1;

alta_slice led_r(
	.A(\Equal0~4_combout ),
	.B(\Equal0~5_combout ),
	.C(vcc),
	.D(\Equal0~7_combout ),
	.Cin(),
	.Qin(\led_r~q ),
	.Clk(\clk~inputclkctrl_outclk_X24_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X24_Y18_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\led_r~0_combout ),
	.Cout(),
	.Q(\led_r~q ));
defparam led_r.coord_x = 1;
defparam led_r.coord_y = 11;
defparam led_r.coord_z = 11;
defparam led_r.mask = 16'h78F0;
defparam led_r.modeMux = 1'b0;
defparam led_r.FeedbackMux = 1'b1;
defparam led_r.ShiftMux = 1'b0;
defparam led_r.BypassEn = 1'b0;
defparam led_r.CarryEnb = 1'b1;

alta_dio \led~output (
	.padio(led),
	.datain(\led_r~q ),
	.datainh(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \led~output .coord_x = 0;
defparam \led~output .coord_y = 15;
defparam \led~output .coord_z = 2;
defparam \led~output .IN_ASYNC_MODE = 1'b0;
defparam \led~output .IN_SYNC_MODE = 1'b0;
defparam \led~output .IN_POWERUP = 1'b0;
defparam \led~output .IN_ASYNC_DISABLE = 1'b0;
defparam \led~output .IN_SYNC_DISABLE = 1'b0;
defparam \led~output .OUT_REG_MODE = 1'b0;
defparam \led~output .OUT_ASYNC_MODE = 1'b0;
defparam \led~output .OUT_SYNC_MODE = 1'b0;
defparam \led~output .OUT_POWERUP = 1'b0;
defparam \led~output .OUT_CLKEN_DISABLE = 1'b0;
defparam \led~output .OUT_ASYNC_DISABLE = 1'b0;
defparam \led~output .OUT_SYNC_DISABLE = 1'b0;
defparam \led~output .OUT_DDIO = 1'b0;
defparam \led~output .OE_REG_MODE = 1'b0;
defparam \led~output .OE_ASYNC_MODE = 1'b0;
defparam \led~output .OE_SYNC_MODE = 1'b0;
defparam \led~output .OE_POWERUP = 1'b0;
defparam \led~output .OE_CLKEN_DISABLE = 1'b0;
defparam \led~output .OE_ASYNC_DISABLE = 1'b0;
defparam \led~output .OE_SYNC_DISABLE = 1'b0;
defparam \led~output .OE_DDIO = 1'b0;
defparam \led~output .CFG_TRI_INPUT = 1'b0;
defparam \led~output .CFG_PULL_UP = 1'b0;
defparam \led~output .CFG_OPEN_DRAIN = 1'b0;
defparam \led~output .CFG_ROCT_CAL_EN = 1'b0;
defparam \led~output .CFG_PDRV = 7'b0011010;
defparam \led~output .CFG_NDRV = 7'b0011000;
defparam \led~output .CFG_KEEP = 2'b00;
defparam \led~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \led~output .CFG_LVDS_SEL_CUA = 3'b000;
defparam \led~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \led~output .CFG_LVDS_IN_EN = 1'b0;
defparam \led~output .CFG_SSTL_OUT_EN = 1'b0;
defparam \led~output .CFG_SSTL_INPUT_EN = 1'b0;
defparam \led~output .CFG_SSTL_SEL_CUA = 3'b011;
defparam \led~output .CFG_OSCDIV = 2'b00;
defparam \led~output .CFG_ROCTUSR = 1'b0;
defparam \led~output .CFG_SEL_CUA = 1'b0;
defparam \led~output .CFG_ROCT_EN = 1'b0;
defparam \led~output .INPUT_ONLY = 1'b0;
defparam \led~output .DPCLK_DELAY = 4'b0000;
defparam \led~output .OUT_DELAY = 1'b0;
defparam \led~output .IN_DATA_DELAY = 3'b000;
defparam \led~output .IN_REG_DELAY = 3'b000;

alta_slice \mii_to_rmii_inst|eth_tx_data[0] (
	.A(\mii_to_rmii_inst|eth_tx_data_reg [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\mii_to_rmii_inst|eth_tx_data [0]),
	.Clk(\e_rxclk~input_o_X33_Y16_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|eth_tx_data[0]~feeder_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|eth_tx_data [0]));
defparam \mii_to_rmii_inst|eth_tx_data[0] .coord_x = 24;
defparam \mii_to_rmii_inst|eth_tx_data[0] .coord_y = 9;
defparam \mii_to_rmii_inst|eth_tx_data[0] .coord_z = 13;
defparam \mii_to_rmii_inst|eth_tx_data[0] .mask = 16'hAAAA;
defparam \mii_to_rmii_inst|eth_tx_data[0] .modeMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[0] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[0] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[0] .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[0] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|eth_tx_data[1] (
	.A(vcc),
	.B(\mii_to_rmii_inst|eth_tx_data_reg [1]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\mii_to_rmii_inst|eth_tx_data [1]),
	.Clk(\e_rxclk~input_o_X33_Y16_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|eth_tx_data[1]~feeder_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|eth_tx_data [1]));
defparam \mii_to_rmii_inst|eth_tx_data[1] .coord_x = 24;
defparam \mii_to_rmii_inst|eth_tx_data[1] .coord_y = 9;
defparam \mii_to_rmii_inst|eth_tx_data[1] .coord_z = 2;
defparam \mii_to_rmii_inst|eth_tx_data[1] .mask = 16'hCCCC;
defparam \mii_to_rmii_inst|eth_tx_data[1] .modeMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[1] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[1] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[1] .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data[1] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|eth_tx_data_reg[0] (
	.A(\mii_to_rmii_inst|tx_data_reg [2]),
	.B(\mii_to_rmii_inst|tx_data_reg [0]),
	.C(vcc),
	.D(\mii_to_rmii_inst|rd_flag~q ),
	.Cin(),
	.Qin(\mii_to_rmii_inst|eth_tx_data_reg [0]),
	.Clk(\e_rxclk~input_o__mii_to_rmii_inst|tx_dv_reg~q_X33_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|eth_tx_data_reg~0_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|eth_tx_data_reg [0]));
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .coord_x = 24;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .coord_y = 9;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .coord_z = 15;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .mask = 16'hAACC;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .modeMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[0] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|eth_tx_data_reg[1] (
	.A(vcc),
	.B(\mii_to_rmii_inst|tx_data_reg [3]),
	.C(\mii_to_rmii_inst|tx_data_reg [1]),
	.D(\mii_to_rmii_inst|rd_flag~q ),
	.Cin(),
	.Qin(\mii_to_rmii_inst|eth_tx_data_reg [1]),
	.Clk(\e_rxclk~input_o__mii_to_rmii_inst|tx_dv_reg~q_X33_Y16_SIG_SIG ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|eth_tx_data_reg~1_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|eth_tx_data_reg [1]));
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .coord_x = 24;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .coord_y = 9;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .coord_z = 7;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .mask = 16'hCCF0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .modeMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_data_reg[1] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|eth_tx_dv (
	.A(\mii_to_rmii_inst|tx_dv_reg~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\mii_to_rmii_inst|eth_tx_dv~q ),
	.Clk(\e_rxclk~input_o_X33_Y16_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|eth_tx_dv~feeder_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|eth_tx_dv~q ));
defparam \mii_to_rmii_inst|eth_tx_dv .coord_x = 24;
defparam \mii_to_rmii_inst|eth_tx_dv .coord_y = 9;
defparam \mii_to_rmii_inst|eth_tx_dv .coord_z = 0;
defparam \mii_to_rmii_inst|eth_tx_dv .mask = 16'hAAAA;
defparam \mii_to_rmii_inst|eth_tx_dv .modeMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_dv .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_dv .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_dv .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|eth_tx_dv .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|rd_flag (
	.A(\mii_to_rmii_inst|tx_dv_reg~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\mii_to_rmii_inst|rd_flag~q ),
	.Clk(\e_rxclk~input_o_X33_Y16_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|rd_flag~0_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|rd_flag~q ));
defparam \mii_to_rmii_inst|rd_flag .coord_x = 24;
defparam \mii_to_rmii_inst|rd_flag .coord_y = 9;
defparam \mii_to_rmii_inst|rd_flag .coord_z = 3;
defparam \mii_to_rmii_inst|rd_flag .mask = 16'h0A0A;
defparam \mii_to_rmii_inst|rd_flag .modeMux = 1'b0;
defparam \mii_to_rmii_inst|rd_flag .FeedbackMux = 1'b1;
defparam \mii_to_rmii_inst|rd_flag .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|rd_flag .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|rd_flag .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|tx_data_reg[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [0]),
	.Cin(),
	.Qin(\mii_to_rmii_inst|tx_data_reg [0]),
	.Clk(\e_rxclk~input_o_X33_Y16_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|tx_data_reg[0]~feeder_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|tx_data_reg [0]));
defparam \mii_to_rmii_inst|tx_data_reg[0] .coord_x = 24;
defparam \mii_to_rmii_inst|tx_data_reg[0] .coord_y = 9;
defparam \mii_to_rmii_inst|tx_data_reg[0] .coord_z = 10;
defparam \mii_to_rmii_inst|tx_data_reg[0] .mask = 16'hFF00;
defparam \mii_to_rmii_inst|tx_data_reg[0] .modeMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[0] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[0] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[0] .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[0] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|tx_data_reg[1] (
	.A(),
	.B(),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [1]),
	.D(),
	.Cin(),
	.Qin(\mii_to_rmii_inst|tx_data_reg [1]),
	.Clk(\e_rxclk~input_o_X33_Y16_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ),
	.SyncReset(SyncReset_X33_Y16_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X33_Y16_VCC),
	.LutOut(),
	.Cout(),
	.Q(\mii_to_rmii_inst|tx_data_reg [1]));
defparam \mii_to_rmii_inst|tx_data_reg[1] .coord_x = 24;
defparam \mii_to_rmii_inst|tx_data_reg[1] .coord_y = 9;
defparam \mii_to_rmii_inst|tx_data_reg[1] .coord_z = 14;
defparam \mii_to_rmii_inst|tx_data_reg[1] .mask = 16'hFFFF;
defparam \mii_to_rmii_inst|tx_data_reg[1] .modeMux = 1'b1;
defparam \mii_to_rmii_inst|tx_data_reg[1] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[1] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[1] .BypassEn = 1'b1;
defparam \mii_to_rmii_inst|tx_data_reg[1] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|tx_data_reg[2] (
	.A(vcc),
	.B(vcc),
	.C(\eth_udp_inst|ip_send_inst|eth_tx_data [2]),
	.D(vcc),
	.Cin(),
	.Qin(\mii_to_rmii_inst|tx_data_reg [2]),
	.Clk(\e_rxclk~input_o_X33_Y16_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|tx_data_reg[2]~feeder_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|tx_data_reg [2]));
defparam \mii_to_rmii_inst|tx_data_reg[2] .coord_x = 24;
defparam \mii_to_rmii_inst|tx_data_reg[2] .coord_y = 9;
defparam \mii_to_rmii_inst|tx_data_reg[2] .coord_z = 5;
defparam \mii_to_rmii_inst|tx_data_reg[2] .mask = 16'hF0F0;
defparam \mii_to_rmii_inst|tx_data_reg[2] .modeMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[2] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[2] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[2] .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[2] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|tx_data_reg[3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_data [3]),
	.Cin(),
	.Qin(\mii_to_rmii_inst|tx_data_reg [3]),
	.Clk(\e_rxclk~input_o_X33_Y16_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|tx_data_reg[3]~feeder_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|tx_data_reg [3]));
defparam \mii_to_rmii_inst|tx_data_reg[3] .coord_x = 24;
defparam \mii_to_rmii_inst|tx_data_reg[3] .coord_y = 9;
defparam \mii_to_rmii_inst|tx_data_reg[3] .coord_z = 8;
defparam \mii_to_rmii_inst|tx_data_reg[3] .mask = 16'hFF00;
defparam \mii_to_rmii_inst|tx_data_reg[3] .modeMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[3] .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[3] .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[3] .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|tx_data_reg[3] .CarryEnb = 1'b1;

alta_slice \mii_to_rmii_inst|tx_dv_reg (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\eth_udp_inst|ip_send_inst|eth_tx_en~q ),
	.Cin(),
	.Qin(\mii_to_rmii_inst|tx_dv_reg~q ),
	.Clk(\e_rxclk~input_o_X33_Y16_INV_VCC ),
	.AsyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~clkctrl_outclk__AsyncReset_X33_Y16_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\mii_to_rmii_inst|tx_dv_reg~feeder_combout ),
	.Cout(),
	.Q(\mii_to_rmii_inst|tx_dv_reg~q ));
defparam \mii_to_rmii_inst|tx_dv_reg .coord_x = 24;
defparam \mii_to_rmii_inst|tx_dv_reg .coord_y = 9;
defparam \mii_to_rmii_inst|tx_dv_reg .coord_z = 11;
defparam \mii_to_rmii_inst|tx_dv_reg .mask = 16'hFF00;
defparam \mii_to_rmii_inst|tx_dv_reg .modeMux = 1'b0;
defparam \mii_to_rmii_inst|tx_dv_reg .FeedbackMux = 1'b0;
defparam \mii_to_rmii_inst|tx_dv_reg .ShiftMux = 1'b0;
defparam \mii_to_rmii_inst|tx_dv_reg .BypassEn = 1'b0;
defparam \mii_to_rmii_inst|tx_dv_reg .CarryEnb = 1'b1;

alta_slice \reset_init[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(reset_init[0]),
	.Clk(\clk~inputclkctrl_outclk__reset_init[5]_X33_Y12_SIG_INV ),
	.AsyncReset(AsyncReset_X33_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\reset_init[0]~1_combout ),
	.Cout(),
	.Q(reset_init[0]));
defparam \reset_init[0] .coord_x = 47;
defparam \reset_init[0] .coord_y = 15;
defparam \reset_init[0] .coord_z = 13;
defparam \reset_init[0] .mask = 16'h0F0F;
defparam \reset_init[0] .modeMux = 1'b0;
defparam \reset_init[0] .FeedbackMux = 1'b1;
defparam \reset_init[0] .ShiftMux = 1'b0;
defparam \reset_init[0] .BypassEn = 1'b0;
defparam \reset_init[0] .CarryEnb = 1'b1;

alta_slice \reset_init[1] (
	.A(reset_init[0]),
	.B(reset_init[1]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(reset_init[1]),
	.Clk(\clk~inputclkctrl_outclk__reset_init[5]_X33_Y12_SIG_INV ),
	.AsyncReset(AsyncReset_X33_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Add0~0_combout ),
	.Cout(\Add0~1 ),
	.Q(reset_init[1]));
defparam \reset_init[1] .coord_x = 47;
defparam \reset_init[1] .coord_y = 15;
defparam \reset_init[1] .coord_z = 5;
defparam \reset_init[1] .mask = 16'h6688;
defparam \reset_init[1] .modeMux = 1'b0;
defparam \reset_init[1] .FeedbackMux = 1'b0;
defparam \reset_init[1] .ShiftMux = 1'b0;
defparam \reset_init[1] .BypassEn = 1'b0;
defparam \reset_init[1] .CarryEnb = 1'b0;

alta_slice \reset_init[2] (
	.A(reset_init[2]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\Add0~1 ),
	.Qin(reset_init[2]),
	.Clk(\clk~inputclkctrl_outclk__reset_init[5]_X33_Y12_SIG_INV ),
	.AsyncReset(AsyncReset_X33_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Add0~2_combout ),
	.Cout(\Add0~3 ),
	.Q(reset_init[2]));
defparam \reset_init[2] .coord_x = 47;
defparam \reset_init[2] .coord_y = 15;
defparam \reset_init[2] .coord_z = 6;
defparam \reset_init[2] .mask = 16'h5A5F;
defparam \reset_init[2] .modeMux = 1'b1;
defparam \reset_init[2] .FeedbackMux = 1'b0;
defparam \reset_init[2] .ShiftMux = 1'b0;
defparam \reset_init[2] .BypassEn = 1'b0;
defparam \reset_init[2] .CarryEnb = 1'b0;

alta_slice \reset_init[3] (
	.A(vcc),
	.B(reset_init[3]),
	.C(vcc),
	.D(vcc),
	.Cin(\Add0~3 ),
	.Qin(reset_init[3]),
	.Clk(\clk~inputclkctrl_outclk__reset_init[5]_X33_Y12_SIG_INV ),
	.AsyncReset(AsyncReset_X33_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Add0~4_combout ),
	.Cout(\Add0~5 ),
	.Q(reset_init[3]));
defparam \reset_init[3] .coord_x = 47;
defparam \reset_init[3] .coord_y = 15;
defparam \reset_init[3] .coord_z = 7;
defparam \reset_init[3] .mask = 16'hC30C;
defparam \reset_init[3] .modeMux = 1'b1;
defparam \reset_init[3] .FeedbackMux = 1'b0;
defparam \reset_init[3] .ShiftMux = 1'b0;
defparam \reset_init[3] .BypassEn = 1'b0;
defparam \reset_init[3] .CarryEnb = 1'b0;

alta_slice \reset_init[4] (
	.A(vcc),
	.B(reset_init[4]),
	.C(vcc),
	.D(vcc),
	.Cin(\Add0~5 ),
	.Qin(reset_init[4]),
	.Clk(\clk~inputclkctrl_outclk__reset_init[5]_X33_Y12_SIG_INV ),
	.AsyncReset(AsyncReset_X33_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\Add0~6_combout ),
	.Cout(\Add0~7 ),
	.Q(reset_init[4]));
defparam \reset_init[4] .coord_x = 47;
defparam \reset_init[4] .coord_y = 15;
defparam \reset_init[4] .coord_z = 8;
defparam \reset_init[4] .mask = 16'h3C3F;
defparam \reset_init[4] .modeMux = 1'b1;
defparam \reset_init[4] .FeedbackMux = 1'b0;
defparam \reset_init[4] .ShiftMux = 1'b0;
defparam \reset_init[4] .BypassEn = 1'b0;
defparam \reset_init[4] .CarryEnb = 1'b0;

alta_slice \reset_init[5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\Add0~8_combout ),
	.Cin(),
	.Qin(reset_init[5]),
	.Clk(\clk~inputclkctrl_outclk_X33_Y12_SIG_VCC ),
	.AsyncReset(AsyncReset_X33_Y12_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\reset_init[5]~0_combout ),
	.Cout(),
	.Q(reset_init[5]));
defparam \reset_init[5] .coord_x = 47;
defparam \reset_init[5] .coord_y = 15;
defparam \reset_init[5] .coord_z = 4;
defparam \reset_init[5] .mask = 16'hFFF0;
defparam \reset_init[5] .modeMux = 1'b0;
defparam \reset_init[5] .FeedbackMux = 1'b1;
defparam \reset_init[5] .ShiftMux = 1'b0;
defparam \reset_init[5] .BypassEn = 1'b0;
defparam \reset_init[5] .CarryEnb = 1'b1;

alta_io_gclk \reset_init[5]~clkctrl (
	.inclk(reset_init[5]),
	.outclk(\reset_init[5]~clkctrl_outclk ));
defparam \reset_init[5]~clkctrl .coord_x = 49;
defparam \reset_init[5]~clkctrl .coord_y = 15;
defparam \reset_init[5]~clkctrl .coord_z = 3;

alta_dio \rst_n~input (
	.padio(rst_n),
	.datain(gnd),
	.datainh(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\rst_n~input_o ),
	.regout());
defparam \rst_n~input .coord_x = 49;
defparam \rst_n~input .coord_y = 15;
defparam \rst_n~input .coord_z = 0;
defparam \rst_n~input .IN_ASYNC_MODE = 1'b0;
defparam \rst_n~input .IN_SYNC_MODE = 1'b0;
defparam \rst_n~input .IN_POWERUP = 1'b0;
defparam \rst_n~input .IN_ASYNC_DISABLE = 1'b0;
defparam \rst_n~input .IN_SYNC_DISABLE = 1'b0;
defparam \rst_n~input .OUT_REG_MODE = 1'b0;
defparam \rst_n~input .OUT_ASYNC_MODE = 1'b0;
defparam \rst_n~input .OUT_SYNC_MODE = 1'b0;
defparam \rst_n~input .OUT_POWERUP = 1'b0;
defparam \rst_n~input .OUT_CLKEN_DISABLE = 1'b0;
defparam \rst_n~input .OUT_ASYNC_DISABLE = 1'b0;
defparam \rst_n~input .OUT_SYNC_DISABLE = 1'b0;
defparam \rst_n~input .OUT_DDIO = 1'b0;
defparam \rst_n~input .OE_REG_MODE = 1'b0;
defparam \rst_n~input .OE_ASYNC_MODE = 1'b0;
defparam \rst_n~input .OE_SYNC_MODE = 1'b0;
defparam \rst_n~input .OE_POWERUP = 1'b0;
defparam \rst_n~input .OE_CLKEN_DISABLE = 1'b0;
defparam \rst_n~input .OE_ASYNC_DISABLE = 1'b0;
defparam \rst_n~input .OE_SYNC_DISABLE = 1'b0;
defparam \rst_n~input .OE_DDIO = 1'b0;
defparam \rst_n~input .CFG_TRI_INPUT = 1'b0;
defparam \rst_n~input .CFG_PULL_UP = 1'b0;
defparam \rst_n~input .CFG_OPEN_DRAIN = 1'b0;
defparam \rst_n~input .CFG_ROCT_CAL_EN = 1'b0;
defparam \rst_n~input .CFG_PDRV = 7'b0010000;
defparam \rst_n~input .CFG_NDRV = 7'b0010000;
defparam \rst_n~input .CFG_KEEP = 2'b00;
defparam \rst_n~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \rst_n~input .CFG_LVDS_SEL_CUA = 3'b000;
defparam \rst_n~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \rst_n~input .CFG_LVDS_IN_EN = 1'b0;
defparam \rst_n~input .CFG_SSTL_OUT_EN = 1'b0;
defparam \rst_n~input .CFG_SSTL_INPUT_EN = 1'b0;
defparam \rst_n~input .CFG_SSTL_SEL_CUA = 3'b011;
defparam \rst_n~input .CFG_OSCDIV = 2'b00;
defparam \rst_n~input .CFG_ROCTUSR = 1'b0;
defparam \rst_n~input .CFG_SEL_CUA = 1'b0;
defparam \rst_n~input .CFG_ROCT_EN = 1'b0;
defparam \rst_n~input .INPUT_ONLY = 1'b1;
defparam \rst_n~input .DPCLK_DELAY = 4'b0000;
defparam \rst_n~input .OUT_DELAY = 1'b0;
defparam \rst_n~input .IN_DATA_DELAY = 3'b000;
defparam \rst_n~input .IN_REG_DELAY = 3'b000;

alta_syncctrl syncload_ctrl_X10_Y9(
	.Din(),
	.Dout(SyncLoad_X10_Y9_VCC));
defparam syncload_ctrl_X10_Y9.coord_x = 16;
defparam syncload_ctrl_X10_Y9.coord_y = 13;
defparam syncload_ctrl_X10_Y9.coord_z = 1;
defparam syncload_ctrl_X10_Y9.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X11_Y14(
	.Din(),
	.Dout(SyncLoad_X11_Y14_VCC));
defparam syncload_ctrl_X11_Y14.coord_x = 9;
defparam syncload_ctrl_X11_Y14.coord_y = 14;
defparam syncload_ctrl_X11_Y14.coord_z = 1;
defparam syncload_ctrl_X11_Y14.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X11_Y16(
	.Din(),
	.Dout(SyncLoad_X11_Y16_VCC));
defparam syncload_ctrl_X11_Y16.coord_x = 16;
defparam syncload_ctrl_X11_Y16.coord_y = 15;
defparam syncload_ctrl_X11_Y16.coord_z = 1;
defparam syncload_ctrl_X11_Y16.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X11_Y9(
	.Din(),
	.Dout(SyncLoad_X11_Y9_VCC));
defparam syncload_ctrl_X11_Y9.coord_x = 16;
defparam syncload_ctrl_X11_Y9.coord_y = 12;
defparam syncload_ctrl_X11_Y9.coord_z = 1;
defparam syncload_ctrl_X11_Y9.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X12_Y14(
	.Din(),
	.Dout(SyncLoad_X12_Y14_VCC));
defparam syncload_ctrl_X12_Y14.coord_x = 10;
defparam syncload_ctrl_X12_Y14.coord_y = 14;
defparam syncload_ctrl_X12_Y14.coord_z = 1;
defparam syncload_ctrl_X12_Y14.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X12_Y16(
	.Din(),
	.Dout(SyncLoad_X12_Y16_VCC));
defparam syncload_ctrl_X12_Y16.coord_x = 17;
defparam syncload_ctrl_X12_Y16.coord_y = 15;
defparam syncload_ctrl_X12_Y16.coord_z = 1;
defparam syncload_ctrl_X12_Y16.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X12_Y18(
	.Din(),
	.Dout(SyncLoad_X12_Y18_VCC));
defparam syncload_ctrl_X12_Y18.coord_x = 11;
defparam syncload_ctrl_X12_Y18.coord_y = 14;
defparam syncload_ctrl_X12_Y18.coord_z = 1;
defparam syncload_ctrl_X12_Y18.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X13_Y10(
	.Din(),
	.Dout(SyncLoad_X13_Y10_VCC));
defparam syncload_ctrl_X13_Y10.coord_x = 17;
defparam syncload_ctrl_X13_Y10.coord_y = 12;
defparam syncload_ctrl_X13_Y10.coord_z = 1;
defparam syncload_ctrl_X13_Y10.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X13_Y16(
	.Din(),
	.Dout(SyncLoad_X13_Y16_VCC));
defparam syncload_ctrl_X13_Y16.coord_x = 17;
defparam syncload_ctrl_X13_Y16.coord_y = 14;
defparam syncload_ctrl_X13_Y16.coord_z = 1;
defparam syncload_ctrl_X13_Y16.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X13_Y18(
	.Din(),
	.Dout(SyncLoad_X13_Y18_VCC));
defparam syncload_ctrl_X13_Y18.coord_x = 10;
defparam syncload_ctrl_X13_Y18.coord_y = 12;
defparam syncload_ctrl_X13_Y18.coord_z = 1;
defparam syncload_ctrl_X13_Y18.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X13_Y7(
	.Din(),
	.Dout(SyncLoad_X13_Y7_VCC));
defparam syncload_ctrl_X13_Y7.coord_x = 17;
defparam syncload_ctrl_X13_Y7.coord_y = 13;
defparam syncload_ctrl_X13_Y7.coord_z = 1;
defparam syncload_ctrl_X13_Y7.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X14_Y10(
	.Din(),
	.Dout(SyncLoad_X14_Y10_VCC));
defparam syncload_ctrl_X14_Y10.coord_x = 16;
defparam syncload_ctrl_X14_Y10.coord_y = 9;
defparam syncload_ctrl_X14_Y10.coord_z = 1;
defparam syncload_ctrl_X14_Y10.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X14_Y16(
	.Din(),
	.Dout(SyncLoad_X14_Y16_VCC));
defparam syncload_ctrl_X14_Y16.coord_x = 13;
defparam syncload_ctrl_X14_Y16.coord_y = 14;
defparam syncload_ctrl_X14_Y16.coord_z = 1;
defparam syncload_ctrl_X14_Y16.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X14_Y18(
	.Din(),
	.Dout(SyncLoad_X14_Y18_VCC));
defparam syncload_ctrl_X14_Y18.coord_x = 13;
defparam syncload_ctrl_X14_Y18.coord_y = 12;
defparam syncload_ctrl_X14_Y18.coord_z = 1;
defparam syncload_ctrl_X14_Y18.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X14_Y19(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y19_SIG ));
defparam syncload_ctrl_X14_Y19.coord_x = 8;
defparam syncload_ctrl_X14_Y19.coord_y = 9;
defparam syncload_ctrl_X14_Y19.coord_z = 1;
defparam syncload_ctrl_X14_Y19.SyncCtrlMux = 2'b10;

alta_syncctrl syncload_ctrl_X14_Y20(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~1_combout__SyncLoad_X14_Y20_SIG ));
defparam syncload_ctrl_X14_Y20.coord_x = 8;
defparam syncload_ctrl_X14_Y20.coord_y = 10;
defparam syncload_ctrl_X14_Y20.coord_z = 1;
defparam syncload_ctrl_X14_Y20.SyncCtrlMux = 2'b10;

alta_syncctrl syncload_ctrl_X14_Y8(
	.Din(),
	.Dout(SyncLoad_X14_Y8_VCC));
defparam syncload_ctrl_X14_Y8.coord_x = 16;
defparam syncload_ctrl_X14_Y8.coord_y = 10;
defparam syncload_ctrl_X14_Y8.coord_z = 1;
defparam syncload_ctrl_X14_Y8.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X14_Y9(
	.Din(),
	.Dout(SyncLoad_X14_Y9_VCC));
defparam syncload_ctrl_X14_Y9.coord_x = 17;
defparam syncload_ctrl_X14_Y9.coord_y = 11;
defparam syncload_ctrl_X14_Y9.coord_z = 1;
defparam syncload_ctrl_X14_Y9.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X16_Y14(
	.Din(),
	.Dout(SyncLoad_X16_Y14_VCC));
defparam syncload_ctrl_X16_Y14.coord_x = 13;
defparam syncload_ctrl_X16_Y14.coord_y = 15;
defparam syncload_ctrl_X16_Y14.coord_z = 1;
defparam syncload_ctrl_X16_Y14.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X16_Y16(
	.Din(),
	.Dout(SyncLoad_X16_Y16_VCC));
defparam syncload_ctrl_X16_Y16.coord_x = 15;
defparam syncload_ctrl_X16_Y16.coord_y = 15;
defparam syncload_ctrl_X16_Y16.coord_z = 1;
defparam syncload_ctrl_X16_Y16.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X16_Y17(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~combout ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|acq_buf_read_reset~combout__SyncLoad_X16_Y17_SIG ));
defparam syncload_ctrl_X16_Y17.coord_x = 17;
defparam syncload_ctrl_X16_Y17.coord_y = 16;
defparam syncload_ctrl_X16_Y17.coord_z = 1;
defparam syncload_ctrl_X16_Y17.SyncCtrlMux = 2'b10;

alta_syncctrl syncload_ctrl_X16_Y18(
	.Din(),
	.Dout(SyncLoad_X16_Y18_VCC));
defparam syncload_ctrl_X16_Y18.coord_x = 14;
defparam syncload_ctrl_X16_Y18.coord_y = 14;
defparam syncload_ctrl_X16_Y18.coord_z = 1;
defparam syncload_ctrl_X16_Y18.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X16_Y19(
	.Din(),
	.Dout(SyncLoad_X16_Y19_VCC));
defparam syncload_ctrl_X16_Y19.coord_x = 14;
defparam syncload_ctrl_X16_Y19.coord_y = 12;
defparam syncload_ctrl_X16_Y19.coord_z = 1;
defparam syncload_ctrl_X16_Y19.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X16_Y9(
	.Din(),
	.Dout(SyncLoad_X16_Y9_VCC));
defparam syncload_ctrl_X16_Y9.coord_x = 17;
defparam syncload_ctrl_X16_Y9.coord_y = 9;
defparam syncload_ctrl_X16_Y9.coord_z = 1;
defparam syncload_ctrl_X16_Y9.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X17_Y15(
	.Din(),
	.Dout(SyncLoad_X17_Y15_GND));
defparam syncload_ctrl_X17_Y15.coord_x = 5;
defparam syncload_ctrl_X17_Y15.coord_y = 15;
defparam syncload_ctrl_X17_Y15.coord_z = 1;
defparam syncload_ctrl_X17_Y15.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X17_Y16(
	.Din(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.Dout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout__SyncLoad_X17_Y16_SIG ));
defparam syncload_ctrl_X17_Y16.coord_x = 7;
defparam syncload_ctrl_X17_Y16.coord_y = 17;
defparam syncload_ctrl_X17_Y16.coord_z = 1;
defparam syncload_ctrl_X17_Y16.SyncCtrlMux = 2'b10;

alta_syncctrl syncload_ctrl_X17_Y17(
	.Din(),
	.Dout(SyncLoad_X17_Y17_VCC));
defparam syncload_ctrl_X17_Y17.coord_x = 6;
defparam syncload_ctrl_X17_Y17.coord_y = 16;
defparam syncload_ctrl_X17_Y17.coord_z = 1;
defparam syncload_ctrl_X17_Y17.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X17_Y20(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0_combout ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_advance_pointer_counter|auto_generated|counter_reg_bit[3]~0_combout__SyncLoad_X17_Y20_SIG ));
defparam syncload_ctrl_X17_Y20.coord_x = 14;
defparam syncload_ctrl_X17_Y20.coord_y = 16;
defparam syncload_ctrl_X17_Y20.coord_z = 1;
defparam syncload_ctrl_X17_Y20.SyncCtrlMux = 2'b10;

alta_syncctrl syncload_ctrl_X17_Y9(
	.Din(),
	.Dout(SyncLoad_X17_Y9_VCC));
defparam syncload_ctrl_X17_Y9.coord_x = 15;
defparam syncload_ctrl_X17_Y9.coord_y = 9;
defparam syncload_ctrl_X17_Y9.coord_z = 1;
defparam syncload_ctrl_X17_Y9.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X18_Y13(
	.Din(),
	.Dout(SyncLoad_X18_Y13_GND));
defparam syncload_ctrl_X18_Y13.coord_x = 5;
defparam syncload_ctrl_X18_Y13.coord_y = 17;
defparam syncload_ctrl_X18_Y13.coord_z = 1;
defparam syncload_ctrl_X18_Y13.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X18_Y15(
	.Din(),
	.Dout(SyncLoad_X18_Y15_GND));
defparam syncload_ctrl_X18_Y15.coord_x = 6;
defparam syncload_ctrl_X18_Y15.coord_y = 15;
defparam syncload_ctrl_X18_Y15.coord_z = 1;
defparam syncload_ctrl_X18_Y15.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X18_Y16(
	.Din(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.Dout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout__SyncLoad_X18_Y16_SIG ));
defparam syncload_ctrl_X18_Y16.coord_x = 6;
defparam syncload_ctrl_X18_Y16.coord_y = 17;
defparam syncload_ctrl_X18_Y16.coord_z = 1;
defparam syncload_ctrl_X18_Y16.SyncCtrlMux = 2'b10;

alta_syncctrl syncload_ctrl_X18_Y17(
	.Din(),
	.Dout(SyncLoad_X18_Y17_VCC));
defparam syncload_ctrl_X18_Y17.coord_x = 5;
defparam syncload_ctrl_X18_Y17.coord_y = 16;
defparam syncload_ctrl_X18_Y17.coord_z = 1;
defparam syncload_ctrl_X18_Y17.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X18_Y18(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena~combout ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|offload_shift_ena~combout__SyncLoad_X18_Y18_INV ));
defparam syncload_ctrl_X18_Y18.coord_x = 8;
defparam syncload_ctrl_X18_Y18.coord_y = 16;
defparam syncload_ctrl_X18_Y18.coord_z = 1;
defparam syncload_ctrl_X18_Y18.SyncCtrlMux = 2'b11;

alta_syncctrl syncload_ctrl_X18_Y19(
	.Din(),
	.Dout(SyncLoad_X18_Y19_VCC));
defparam syncload_ctrl_X18_Y19.coord_x = 10;
defparam syncload_ctrl_X18_Y19.coord_y = 15;
defparam syncload_ctrl_X18_Y19.coord_z = 1;
defparam syncload_ctrl_X18_Y19.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X18_Y20(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0_combout ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|stp_non_zero_depth_offload_gen:stp_offload_buff_mgr_inst|status_read_pointer_counter|auto_generated|counter_reg_bit[0]~0_combout__SyncLoad_X18_Y20_SIG ));
defparam syncload_ctrl_X18_Y20.coord_x = 13;
defparam syncload_ctrl_X18_Y20.coord_y = 16;
defparam syncload_ctrl_X18_Y20.coord_z = 1;
defparam syncload_ctrl_X18_Y20.SyncCtrlMux = 2'b10;

alta_syncctrl syncload_ctrl_X19_Y16(
	.Din(),
	.Dout(SyncLoad_X19_Y16_VCC));
defparam syncload_ctrl_X19_Y16.coord_x = 4;
defparam syncload_ctrl_X19_Y16.coord_y = 17;
defparam syncload_ctrl_X19_Y16.coord_z = 1;
defparam syncload_ctrl_X19_Y16.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X19_Y17(
	.Din(),
	.Dout(SyncLoad_X19_Y17_VCC));
defparam syncload_ctrl_X19_Y17.coord_x = 2;
defparam syncload_ctrl_X19_Y17.coord_y = 15;
defparam syncload_ctrl_X19_Y17.coord_z = 1;
defparam syncload_ctrl_X19_Y17.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X19_Y8(
	.Din(),
	.Dout(SyncLoad_X19_Y8_GND));
defparam syncload_ctrl_X19_Y8.coord_x = 26;
defparam syncload_ctrl_X19_Y8.coord_y = 6;
defparam syncload_ctrl_X19_Y8.coord_z = 1;
defparam syncload_ctrl_X19_Y8.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X1_Y7(
	.Din(),
	.Dout(SyncLoad_X1_Y7_GND));
defparam syncload_ctrl_X1_Y7.coord_x = 4;
defparam syncload_ctrl_X1_Y7.coord_y = 11;
defparam syncload_ctrl_X1_Y7.coord_z = 1;
defparam syncload_ctrl_X1_Y7.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X21_Y15(
	.Din(),
	.Dout(SyncLoad_X21_Y15_GND));
defparam syncload_ctrl_X21_Y15.coord_x = 3;
defparam syncload_ctrl_X21_Y15.coord_y = 15;
defparam syncload_ctrl_X21_Y15.coord_z = 1;
defparam syncload_ctrl_X21_Y15.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X21_Y16(
	.Din(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.Dout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3]__SyncLoad_X21_Y16_SIG ));
defparam syncload_ctrl_X21_Y16.coord_x = 4;
defparam syncload_ctrl_X21_Y16.coord_y = 15;
defparam syncload_ctrl_X21_Y16.coord_z = 1;
defparam syncload_ctrl_X21_Y16.SyncCtrlMux = 2'b10;

alta_syncctrl syncload_ctrl_X21_Y17(
	.Din(),
	.Dout(SyncLoad_X21_Y17_GND));
defparam syncload_ctrl_X21_Y17.coord_x = 1;
defparam syncload_ctrl_X21_Y17.coord_y = 15;
defparam syncload_ctrl_X21_Y17.coord_z = 1;
defparam syncload_ctrl_X21_Y17.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X21_Y18(
	.Din(),
	.Dout(SyncLoad_X21_Y18_VCC));
defparam syncload_ctrl_X21_Y18.coord_x = 9;
defparam syncload_ctrl_X21_Y18.coord_y = 16;
defparam syncload_ctrl_X21_Y18.coord_z = 1;
defparam syncload_ctrl_X21_Y18.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X21_Y19(
	.Din(),
	.Dout(SyncLoad_X21_Y19_VCC));
defparam syncload_ctrl_X21_Y19.coord_x = 11;
defparam syncload_ctrl_X21_Y19.coord_y = 15;
defparam syncload_ctrl_X21_Y19.coord_z = 1;
defparam syncload_ctrl_X21_Y19.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X22_Y14(
	.Din(\eth_udp_inst|ip_send_inst|Equal1~1_combout ),
	.Dout(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y14_SIG ));
defparam syncload_ctrl_X22_Y14.coord_x = 21;
defparam syncload_ctrl_X22_Y14.coord_y = 13;
defparam syncload_ctrl_X22_Y14.coord_z = 1;
defparam syncload_ctrl_X22_Y14.SyncCtrlMux = 2'b10;

alta_syncctrl syncload_ctrl_X22_Y15(
	.Din(\eth_udp_inst|ip_send_inst|Equal1~1_combout ),
	.Dout(\eth_udp_inst|ip_send_inst|Equal1~1_combout__SyncLoad_X22_Y15_SIG ));
defparam syncload_ctrl_X22_Y15.coord_x = 21;
defparam syncload_ctrl_X22_Y15.coord_y = 14;
defparam syncload_ctrl_X22_Y15.coord_z = 1;
defparam syncload_ctrl_X22_Y15.SyncCtrlMux = 2'b10;

alta_syncctrl syncload_ctrl_X23_Y16(
	.Din(),
	.Dout(SyncLoad_X23_Y16_VCC));
defparam syncload_ctrl_X23_Y16.coord_x = 20;
defparam syncload_ctrl_X23_Y16.coord_y = 10;
defparam syncload_ctrl_X23_Y16.coord_z = 1;
defparam syncload_ctrl_X23_Y16.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X24_Y15(
	.Din(),
	.Dout(SyncLoad_X24_Y15_GND));
defparam syncload_ctrl_X24_Y15.coord_x = 21;
defparam syncload_ctrl_X24_Y15.coord_y = 10;
defparam syncload_ctrl_X24_Y15.coord_z = 1;
defparam syncload_ctrl_X24_Y15.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X24_Y16(
	.Din(),
	.Dout(SyncLoad_X24_Y16_VCC));
defparam syncload_ctrl_X24_Y16.coord_x = 20;
defparam syncload_ctrl_X24_Y16.coord_y = 12;
defparam syncload_ctrl_X24_Y16.coord_z = 1;
defparam syncload_ctrl_X24_Y16.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X24_Y19(
	.Din(),
	.Dout(SyncLoad_X24_Y19_VCC));
defparam syncload_ctrl_X24_Y19.coord_x = 12;
defparam syncload_ctrl_X24_Y19.coord_y = 16;
defparam syncload_ctrl_X24_Y19.coord_z = 1;
defparam syncload_ctrl_X24_Y19.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X25_Y12(
	.Din(),
	.Dout(SyncLoad_X25_Y12_VCC));
defparam syncload_ctrl_X25_Y12.coord_x = 21;
defparam syncload_ctrl_X25_Y12.coord_y = 9;
defparam syncload_ctrl_X25_Y12.coord_z = 1;
defparam syncload_ctrl_X25_Y12.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X25_Y18(
	.Din(),
	.Dout(SyncLoad_X25_Y18_GND));
defparam syncload_ctrl_X25_Y18.coord_x = 2;
defparam syncload_ctrl_X25_Y18.coord_y = 11;
defparam syncload_ctrl_X25_Y18.coord_z = 1;
defparam syncload_ctrl_X25_Y18.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X25_Y19(
	.Din(),
	.Dout(SyncLoad_X25_Y19_GND));
defparam syncload_ctrl_X25_Y19.coord_x = 2;
defparam syncload_ctrl_X25_Y19.coord_y = 12;
defparam syncload_ctrl_X25_Y19.coord_z = 1;
defparam syncload_ctrl_X25_Y19.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X26_Y15(
	.Din(),
	.Dout(SyncLoad_X26_Y15_GND));
defparam syncload_ctrl_X26_Y15.coord_x = 19;
defparam syncload_ctrl_X26_Y15.coord_y = 14;
defparam syncload_ctrl_X26_Y15.coord_z = 1;
defparam syncload_ctrl_X26_Y15.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X26_Y16(
	.Din(),
	.Dout(SyncLoad_X26_Y16_GND));
defparam syncload_ctrl_X26_Y16.coord_x = 19;
defparam syncload_ctrl_X26_Y16.coord_y = 12;
defparam syncload_ctrl_X26_Y16.coord_z = 1;
defparam syncload_ctrl_X26_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X28_Y9(
	.Din(),
	.Dout(SyncLoad_X28_Y9_VCC));
defparam syncload_ctrl_X28_Y9.coord_x = 24;
defparam syncload_ctrl_X28_Y9.coord_y = 8;
defparam syncload_ctrl_X28_Y9.coord_z = 1;
defparam syncload_ctrl_X28_Y9.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X29_Y9(
	.Din(),
	.Dout(SyncLoad_X29_Y9_GND));
defparam syncload_ctrl_X29_Y9.coord_x = 25;
defparam syncload_ctrl_X29_Y9.coord_y = 8;
defparam syncload_ctrl_X29_Y9.coord_z = 1;
defparam syncload_ctrl_X29_Y9.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X2_Y7(
	.Din(),
	.Dout(SyncLoad_X2_Y7_VCC));
defparam syncload_ctrl_X2_Y7.coord_x = 5;
defparam syncload_ctrl_X2_Y7.coord_y = 11;
defparam syncload_ctrl_X2_Y7.coord_z = 1;
defparam syncload_ctrl_X2_Y7.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X33_Y16(
	.Din(),
	.Dout(SyncLoad_X33_Y16_VCC));
defparam syncload_ctrl_X33_Y16.coord_x = 24;
defparam syncload_ctrl_X33_Y16.coord_y = 9;
defparam syncload_ctrl_X33_Y16.coord_z = 1;
defparam syncload_ctrl_X33_Y16.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X5_Y7(
	.Din(),
	.Dout(SyncLoad_X5_Y7_GND));
defparam syncload_ctrl_X5_Y7.coord_x = 8;
defparam syncload_ctrl_X5_Y7.coord_y = 11;
defparam syncload_ctrl_X5_Y7.coord_z = 1;
defparam syncload_ctrl_X5_Y7.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X9_Y7(
	.Din(),
	.Dout(SyncLoad_X9_Y7_VCC));
defparam syncload_ctrl_X9_Y7.coord_x = 10;
defparam syncload_ctrl_X9_Y7.coord_y = 11;
defparam syncload_ctrl_X9_Y7.coord_z = 1;
defparam syncload_ctrl_X9_Y7.SyncCtrlMux = 2'b01;

alta_syncctrl syncreset_ctrl_X10_Y9(
	.Din(),
	.Dout(SyncReset_X10_Y9_GND));
defparam syncreset_ctrl_X10_Y9.coord_x = 16;
defparam syncreset_ctrl_X10_Y9.coord_y = 13;
defparam syncreset_ctrl_X10_Y9.coord_z = 0;
defparam syncreset_ctrl_X10_Y9.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X11_Y14(
	.Din(),
	.Dout(SyncReset_X11_Y14_GND));
defparam syncreset_ctrl_X11_Y14.coord_x = 9;
defparam syncreset_ctrl_X11_Y14.coord_y = 14;
defparam syncreset_ctrl_X11_Y14.coord_z = 0;
defparam syncreset_ctrl_X11_Y14.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X11_Y16(
	.Din(),
	.Dout(SyncReset_X11_Y16_GND));
defparam syncreset_ctrl_X11_Y16.coord_x = 16;
defparam syncreset_ctrl_X11_Y16.coord_y = 15;
defparam syncreset_ctrl_X11_Y16.coord_z = 0;
defparam syncreset_ctrl_X11_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X11_Y9(
	.Din(),
	.Dout(SyncReset_X11_Y9_GND));
defparam syncreset_ctrl_X11_Y9.coord_x = 16;
defparam syncreset_ctrl_X11_Y9.coord_y = 12;
defparam syncreset_ctrl_X11_Y9.coord_z = 0;
defparam syncreset_ctrl_X11_Y9.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X12_Y14(
	.Din(),
	.Dout(SyncReset_X12_Y14_GND));
defparam syncreset_ctrl_X12_Y14.coord_x = 10;
defparam syncreset_ctrl_X12_Y14.coord_y = 14;
defparam syncreset_ctrl_X12_Y14.coord_z = 0;
defparam syncreset_ctrl_X12_Y14.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X12_Y16(
	.Din(),
	.Dout(SyncReset_X12_Y16_GND));
defparam syncreset_ctrl_X12_Y16.coord_x = 17;
defparam syncreset_ctrl_X12_Y16.coord_y = 15;
defparam syncreset_ctrl_X12_Y16.coord_z = 0;
defparam syncreset_ctrl_X12_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X12_Y18(
	.Din(),
	.Dout(SyncReset_X12_Y18_GND));
defparam syncreset_ctrl_X12_Y18.coord_x = 11;
defparam syncreset_ctrl_X12_Y18.coord_y = 14;
defparam syncreset_ctrl_X12_Y18.coord_z = 0;
defparam syncreset_ctrl_X12_Y18.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X13_Y10(
	.Din(),
	.Dout(SyncReset_X13_Y10_GND));
defparam syncreset_ctrl_X13_Y10.coord_x = 17;
defparam syncreset_ctrl_X13_Y10.coord_y = 12;
defparam syncreset_ctrl_X13_Y10.coord_z = 0;
defparam syncreset_ctrl_X13_Y10.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X13_Y16(
	.Din(),
	.Dout(SyncReset_X13_Y16_GND));
defparam syncreset_ctrl_X13_Y16.coord_x = 17;
defparam syncreset_ctrl_X13_Y16.coord_y = 14;
defparam syncreset_ctrl_X13_Y16.coord_z = 0;
defparam syncreset_ctrl_X13_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X13_Y18(
	.Din(),
	.Dout(SyncReset_X13_Y18_GND));
defparam syncreset_ctrl_X13_Y18.coord_x = 10;
defparam syncreset_ctrl_X13_Y18.coord_y = 12;
defparam syncreset_ctrl_X13_Y18.coord_z = 0;
defparam syncreset_ctrl_X13_Y18.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X13_Y7(
	.Din(),
	.Dout(SyncReset_X13_Y7_GND));
defparam syncreset_ctrl_X13_Y7.coord_x = 17;
defparam syncreset_ctrl_X13_Y7.coord_y = 13;
defparam syncreset_ctrl_X13_Y7.coord_z = 0;
defparam syncreset_ctrl_X13_Y7.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X14_Y10(
	.Din(),
	.Dout(SyncReset_X14_Y10_GND));
defparam syncreset_ctrl_X14_Y10.coord_x = 16;
defparam syncreset_ctrl_X14_Y10.coord_y = 9;
defparam syncreset_ctrl_X14_Y10.coord_z = 0;
defparam syncreset_ctrl_X14_Y10.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X14_Y16(
	.Din(),
	.Dout(SyncReset_X14_Y16_GND));
defparam syncreset_ctrl_X14_Y16.coord_x = 13;
defparam syncreset_ctrl_X14_Y16.coord_y = 14;
defparam syncreset_ctrl_X14_Y16.coord_z = 0;
defparam syncreset_ctrl_X14_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X14_Y18(
	.Din(),
	.Dout(SyncReset_X14_Y18_GND));
defparam syncreset_ctrl_X14_Y18.coord_x = 13;
defparam syncreset_ctrl_X14_Y18.coord_y = 12;
defparam syncreset_ctrl_X14_Y18.coord_z = 0;
defparam syncreset_ctrl_X14_Y18.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X14_Y19(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y19_SIG ));
defparam syncreset_ctrl_X14_Y19.coord_x = 8;
defparam syncreset_ctrl_X14_Y19.coord_y = 9;
defparam syncreset_ctrl_X14_Y19.coord_z = 0;
defparam syncreset_ctrl_X14_Y19.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X14_Y20(
	.Din(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout ),
	.Dout(\auto_signaltap_0|sld_signaltap_body|sld_signaltap_body|process_0~0_combout__SyncReset_X14_Y20_SIG ));
defparam syncreset_ctrl_X14_Y20.coord_x = 8;
defparam syncreset_ctrl_X14_Y20.coord_y = 10;
defparam syncreset_ctrl_X14_Y20.coord_z = 0;
defparam syncreset_ctrl_X14_Y20.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X14_Y8(
	.Din(),
	.Dout(SyncReset_X14_Y8_GND));
defparam syncreset_ctrl_X14_Y8.coord_x = 16;
defparam syncreset_ctrl_X14_Y8.coord_y = 10;
defparam syncreset_ctrl_X14_Y8.coord_z = 0;
defparam syncreset_ctrl_X14_Y8.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X14_Y9(
	.Din(),
	.Dout(SyncReset_X14_Y9_GND));
defparam syncreset_ctrl_X14_Y9.coord_x = 17;
defparam syncreset_ctrl_X14_Y9.coord_y = 11;
defparam syncreset_ctrl_X14_Y9.coord_z = 0;
defparam syncreset_ctrl_X14_Y9.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X16_Y14(
	.Din(),
	.Dout(SyncReset_X16_Y14_GND));
defparam syncreset_ctrl_X16_Y14.coord_x = 13;
defparam syncreset_ctrl_X16_Y14.coord_y = 15;
defparam syncreset_ctrl_X16_Y14.coord_z = 0;
defparam syncreset_ctrl_X16_Y14.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X16_Y16(
	.Din(),
	.Dout(SyncReset_X16_Y16_GND));
defparam syncreset_ctrl_X16_Y16.coord_x = 15;
defparam syncreset_ctrl_X16_Y16.coord_y = 15;
defparam syncreset_ctrl_X16_Y16.coord_z = 0;
defparam syncreset_ctrl_X16_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X16_Y17(
	.Din(),
	.Dout(SyncReset_X16_Y17_GND));
defparam syncreset_ctrl_X16_Y17.coord_x = 17;
defparam syncreset_ctrl_X16_Y17.coord_y = 16;
defparam syncreset_ctrl_X16_Y17.coord_z = 0;
defparam syncreset_ctrl_X16_Y17.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X16_Y18(
	.Din(),
	.Dout(SyncReset_X16_Y18_GND));
defparam syncreset_ctrl_X16_Y18.coord_x = 14;
defparam syncreset_ctrl_X16_Y18.coord_y = 14;
defparam syncreset_ctrl_X16_Y18.coord_z = 0;
defparam syncreset_ctrl_X16_Y18.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X16_Y19(
	.Din(),
	.Dout(SyncReset_X16_Y19_GND));
defparam syncreset_ctrl_X16_Y19.coord_x = 14;
defparam syncreset_ctrl_X16_Y19.coord_y = 12;
defparam syncreset_ctrl_X16_Y19.coord_z = 0;
defparam syncreset_ctrl_X16_Y19.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X16_Y9(
	.Din(),
	.Dout(SyncReset_X16_Y9_GND));
defparam syncreset_ctrl_X16_Y9.coord_x = 17;
defparam syncreset_ctrl_X16_Y9.coord_y = 9;
defparam syncreset_ctrl_X16_Y9.coord_z = 0;
defparam syncreset_ctrl_X16_Y9.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X17_Y15(
	.Din(\altera_internal_jtag~TMSUTAP ),
	.Dout(\altera_internal_jtag~TMSUTAP__SyncReset_X17_Y15_SIG ));
defparam syncreset_ctrl_X17_Y15.coord_x = 5;
defparam syncreset_ctrl_X17_Y15.coord_y = 15;
defparam syncreset_ctrl_X17_Y15.coord_z = 0;
defparam syncreset_ctrl_X17_Y15.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X17_Y16(
	.Din(),
	.Dout(SyncReset_X17_Y16_GND));
defparam syncreset_ctrl_X17_Y16.coord_x = 7;
defparam syncreset_ctrl_X17_Y16.coord_y = 17;
defparam syncreset_ctrl_X17_Y16.coord_z = 0;
defparam syncreset_ctrl_X17_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X17_Y17(
	.Din(),
	.Dout(SyncReset_X17_Y17_GND));
defparam syncreset_ctrl_X17_Y17.coord_x = 6;
defparam syncreset_ctrl_X17_Y17.coord_y = 16;
defparam syncreset_ctrl_X17_Y17.coord_z = 0;
defparam syncreset_ctrl_X17_Y17.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X17_Y20(
	.Din(),
	.Dout(SyncReset_X17_Y20_GND));
defparam syncreset_ctrl_X17_Y20.coord_x = 14;
defparam syncreset_ctrl_X17_Y20.coord_y = 16;
defparam syncreset_ctrl_X17_Y20.coord_z = 0;
defparam syncreset_ctrl_X17_Y20.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X17_Y9(
	.Din(),
	.Dout(SyncReset_X17_Y9_GND));
defparam syncreset_ctrl_X17_Y9.coord_x = 15;
defparam syncreset_ctrl_X17_Y9.coord_y = 9;
defparam syncreset_ctrl_X17_Y9.coord_z = 0;
defparam syncreset_ctrl_X17_Y9.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X18_Y13(
	.Din(\altera_internal_jtag~TMSUTAP ),
	.Dout(\altera_internal_jtag~TMSUTAP__SyncReset_X18_Y13_SIG ));
defparam syncreset_ctrl_X18_Y13.coord_x = 5;
defparam syncreset_ctrl_X18_Y13.coord_y = 17;
defparam syncreset_ctrl_X18_Y13.coord_z = 0;
defparam syncreset_ctrl_X18_Y13.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X18_Y15(
	.Din(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13_combout ),
	.Dout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~13_combout__SyncReset_X18_Y15_SIG ));
defparam syncreset_ctrl_X18_Y15.coord_x = 6;
defparam syncreset_ctrl_X18_Y15.coord_y = 15;
defparam syncreset_ctrl_X18_Y15.coord_z = 0;
defparam syncreset_ctrl_X18_Y15.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X18_Y16(
	.Din(),
	.Dout(SyncReset_X18_Y16_GND));
defparam syncreset_ctrl_X18_Y16.coord_x = 6;
defparam syncreset_ctrl_X18_Y16.coord_y = 17;
defparam syncreset_ctrl_X18_Y16.coord_z = 0;
defparam syncreset_ctrl_X18_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X18_Y17(
	.Din(),
	.Dout(SyncReset_X18_Y17_GND));
defparam syncreset_ctrl_X18_Y17.coord_x = 5;
defparam syncreset_ctrl_X18_Y17.coord_y = 16;
defparam syncreset_ctrl_X18_Y17.coord_z = 0;
defparam syncreset_ctrl_X18_Y17.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X18_Y18(
	.Din(),
	.Dout(SyncReset_X18_Y18_GND));
defparam syncreset_ctrl_X18_Y18.coord_x = 8;
defparam syncreset_ctrl_X18_Y18.coord_y = 16;
defparam syncreset_ctrl_X18_Y18.coord_z = 0;
defparam syncreset_ctrl_X18_Y18.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X18_Y19(
	.Din(),
	.Dout(SyncReset_X18_Y19_GND));
defparam syncreset_ctrl_X18_Y19.coord_x = 10;
defparam syncreset_ctrl_X18_Y19.coord_y = 15;
defparam syncreset_ctrl_X18_Y19.coord_z = 0;
defparam syncreset_ctrl_X18_Y19.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X18_Y20(
	.Din(),
	.Dout(SyncReset_X18_Y20_GND));
defparam syncreset_ctrl_X18_Y20.coord_x = 13;
defparam syncreset_ctrl_X18_Y20.coord_y = 16;
defparam syncreset_ctrl_X18_Y20.coord_z = 0;
defparam syncreset_ctrl_X18_Y20.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X19_Y16(
	.Din(),
	.Dout(SyncReset_X19_Y16_GND));
defparam syncreset_ctrl_X19_Y16.coord_x = 4;
defparam syncreset_ctrl_X19_Y16.coord_y = 17;
defparam syncreset_ctrl_X19_Y16.coord_z = 0;
defparam syncreset_ctrl_X19_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X19_Y17(
	.Din(),
	.Dout(SyncReset_X19_Y17_GND));
defparam syncreset_ctrl_X19_Y17.coord_x = 2;
defparam syncreset_ctrl_X19_Y17.coord_y = 15;
defparam syncreset_ctrl_X19_Y17.coord_z = 0;
defparam syncreset_ctrl_X19_Y17.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X19_Y8(
	.Din(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout ),
	.Dout(\camera_if_inst|u_I2C_AV_Config|mI2C_GO~0_combout__SyncReset_X19_Y8_INV ));
defparam syncreset_ctrl_X19_Y8.coord_x = 26;
defparam syncreset_ctrl_X19_Y8.coord_y = 6;
defparam syncreset_ctrl_X19_Y8.coord_z = 0;
defparam syncreset_ctrl_X19_Y8.SyncCtrlMux = 2'b11;

alta_syncctrl syncreset_ctrl_X1_Y7(
	.Din(\camera_if_inst|cam_hsync_r [0]),
	.Dout(\camera_if_inst|cam_hsync_r[0]__SyncReset_X1_Y7_INV ));
defparam syncreset_ctrl_X1_Y7.coord_x = 4;
defparam syncreset_ctrl_X1_Y7.coord_y = 11;
defparam syncreset_ctrl_X1_Y7.coord_z = 0;
defparam syncreset_ctrl_X1_Y7.SyncCtrlMux = 2'b11;

alta_syncctrl syncreset_ctrl_X21_Y15(
	.Din(\altera_internal_jtag~TMSUTAP ),
	.Dout(\altera_internal_jtag~TMSUTAP__SyncReset_X21_Y15_INV ));
defparam syncreset_ctrl_X21_Y15.coord_x = 3;
defparam syncreset_ctrl_X21_Y15.coord_y = 15;
defparam syncreset_ctrl_X21_Y15.coord_z = 0;
defparam syncreset_ctrl_X21_Y15.SyncCtrlMux = 2'b11;

alta_syncctrl syncreset_ctrl_X21_Y16(
	.Din(),
	.Dout(SyncReset_X21_Y16_GND));
defparam syncreset_ctrl_X21_Y16.coord_x = 4;
defparam syncreset_ctrl_X21_Y16.coord_y = 15;
defparam syncreset_ctrl_X21_Y16.coord_z = 0;
defparam syncreset_ctrl_X21_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X21_Y17(
	.Din(\altera_internal_jtag~TMSUTAP ),
	.Dout(\altera_internal_jtag~TMSUTAP__SyncReset_X21_Y17_SIG ));
defparam syncreset_ctrl_X21_Y17.coord_x = 1;
defparam syncreset_ctrl_X21_Y17.coord_y = 15;
defparam syncreset_ctrl_X21_Y17.coord_z = 0;
defparam syncreset_ctrl_X21_Y17.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X21_Y18(
	.Din(),
	.Dout(SyncReset_X21_Y18_GND));
defparam syncreset_ctrl_X21_Y18.coord_x = 9;
defparam syncreset_ctrl_X21_Y18.coord_y = 16;
defparam syncreset_ctrl_X21_Y18.coord_z = 0;
defparam syncreset_ctrl_X21_Y18.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X21_Y19(
	.Din(),
	.Dout(SyncReset_X21_Y19_GND));
defparam syncreset_ctrl_X21_Y19.coord_x = 11;
defparam syncreset_ctrl_X21_Y19.coord_y = 15;
defparam syncreset_ctrl_X21_Y19.coord_z = 0;
defparam syncreset_ctrl_X21_Y19.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X22_Y14(
	.Din(),
	.Dout(SyncReset_X22_Y14_GND));
defparam syncreset_ctrl_X22_Y14.coord_x = 21;
defparam syncreset_ctrl_X22_Y14.coord_y = 13;
defparam syncreset_ctrl_X22_Y14.coord_z = 0;
defparam syncreset_ctrl_X22_Y14.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X22_Y15(
	.Din(),
	.Dout(SyncReset_X22_Y15_GND));
defparam syncreset_ctrl_X22_Y15.coord_x = 21;
defparam syncreset_ctrl_X22_Y15.coord_y = 14;
defparam syncreset_ctrl_X22_Y15.coord_z = 0;
defparam syncreset_ctrl_X22_Y15.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X23_Y16(
	.Din(),
	.Dout(SyncReset_X23_Y16_GND));
defparam syncreset_ctrl_X23_Y16.coord_x = 20;
defparam syncreset_ctrl_X23_Y16.coord_y = 10;
defparam syncreset_ctrl_X23_Y16.coord_z = 0;
defparam syncreset_ctrl_X23_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X24_Y15(
	.Din(\eth_udp_inst|ip_send_inst|cnt[4]~11_combout ),
	.Dout(\eth_udp_inst|ip_send_inst|cnt[4]~11_combout__SyncReset_X24_Y15_SIG ));
defparam syncreset_ctrl_X24_Y15.coord_x = 21;
defparam syncreset_ctrl_X24_Y15.coord_y = 10;
defparam syncreset_ctrl_X24_Y15.coord_z = 0;
defparam syncreset_ctrl_X24_Y15.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X24_Y16(
	.Din(),
	.Dout(SyncReset_X24_Y16_GND));
defparam syncreset_ctrl_X24_Y16.coord_x = 20;
defparam syncreset_ctrl_X24_Y16.coord_y = 12;
defparam syncreset_ctrl_X24_Y16.coord_z = 0;
defparam syncreset_ctrl_X24_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X24_Y19(
	.Din(),
	.Dout(SyncReset_X24_Y19_GND));
defparam syncreset_ctrl_X24_Y19.coord_x = 12;
defparam syncreset_ctrl_X24_Y19.coord_y = 16;
defparam syncreset_ctrl_X24_Y19.coord_z = 0;
defparam syncreset_ctrl_X24_Y19.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X25_Y12(
	.Din(),
	.Dout(SyncReset_X25_Y12_GND));
defparam syncreset_ctrl_X25_Y12.coord_x = 21;
defparam syncreset_ctrl_X25_Y12.coord_y = 9;
defparam syncreset_ctrl_X25_Y12.coord_z = 0;
defparam syncreset_ctrl_X25_Y12.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X25_Y18(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ));
defparam syncreset_ctrl_X25_Y18.coord_x = 2;
defparam syncreset_ctrl_X25_Y18.coord_y = 11;
defparam syncreset_ctrl_X25_Y18.coord_z = 0;
defparam syncreset_ctrl_X25_Y18.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X25_Y19(
	.Din(\alt_pll_inst|altpll_component|auto_generated|locked~combout ),
	.Dout(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ));
defparam syncreset_ctrl_X25_Y19.coord_x = 2;
defparam syncreset_ctrl_X25_Y19.coord_y = 12;
defparam syncreset_ctrl_X25_Y19.coord_z = 0;
defparam syncreset_ctrl_X25_Y19.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X26_Y15(
	.Din(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Dout(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y15_SIG ));
defparam syncreset_ctrl_X26_Y15.coord_x = 19;
defparam syncreset_ctrl_X26_Y15.coord_y = 14;
defparam syncreset_ctrl_X26_Y15.coord_z = 0;
defparam syncreset_ctrl_X26_Y15.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X26_Y16(
	.Din(\eth_udp_inst|ip_send_inst|sw_en~q ),
	.Dout(\eth_udp_inst|ip_send_inst|sw_en~q__SyncReset_X26_Y16_SIG ));
defparam syncreset_ctrl_X26_Y16.coord_x = 19;
defparam syncreset_ctrl_X26_Y16.coord_y = 12;
defparam syncreset_ctrl_X26_Y16.coord_z = 0;
defparam syncreset_ctrl_X26_Y16.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X28_Y9(
	.Din(),
	.Dout(SyncReset_X28_Y9_GND));
defparam syncreset_ctrl_X28_Y9.coord_x = 24;
defparam syncreset_ctrl_X28_Y9.coord_y = 8;
defparam syncreset_ctrl_X28_Y9.coord_z = 0;
defparam syncreset_ctrl_X28_Y9.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X29_Y9(
	.Din(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout ),
	.Dout(\camera_if_inst|u_I2C_AV_Config|LessThan0~4_combout__SyncReset_X29_Y9_INV ));
defparam syncreset_ctrl_X29_Y9.coord_x = 25;
defparam syncreset_ctrl_X29_Y9.coord_y = 8;
defparam syncreset_ctrl_X29_Y9.coord_z = 0;
defparam syncreset_ctrl_X29_Y9.SyncCtrlMux = 2'b11;

alta_syncctrl syncreset_ctrl_X2_Y7(
	.Din(),
	.Dout(SyncReset_X2_Y7_GND));
defparam syncreset_ctrl_X2_Y7.coord_x = 5;
defparam syncreset_ctrl_X2_Y7.coord_y = 11;
defparam syncreset_ctrl_X2_Y7.coord_z = 0;
defparam syncreset_ctrl_X2_Y7.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X33_Y16(
	.Din(),
	.Dout(SyncReset_X33_Y16_GND));
defparam syncreset_ctrl_X33_Y16.coord_x = 24;
defparam syncreset_ctrl_X33_Y16.coord_y = 9;
defparam syncreset_ctrl_X33_Y16.coord_z = 0;
defparam syncreset_ctrl_X33_Y16.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X5_Y7(
	.Din(\camera_if_inst|cam_vsync_r [0]),
	.Dout(\camera_if_inst|cam_vsync_r[0]__SyncReset_X5_Y7_SIG ));
defparam syncreset_ctrl_X5_Y7.coord_x = 8;
defparam syncreset_ctrl_X5_Y7.coord_y = 11;
defparam syncreset_ctrl_X5_Y7.coord_z = 0;
defparam syncreset_ctrl_X5_Y7.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X9_Y7(
	.Din(),
	.Dout(SyncReset_X9_Y7_GND));
defparam syncreset_ctrl_X9_Y7.coord_x = 10;
defparam syncreset_ctrl_X9_Y7.coord_y = 11;
defparam syncreset_ctrl_X9_Y7.coord_z = 0;
defparam syncreset_ctrl_X9_Y7.SyncCtrlMux = 2'b00;

alta_slice \timer[0] (
	.A(vcc),
	.B(timer[0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(timer[0]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y19_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y19_GND),
	.LutOut(\timer[0]~25_combout ),
	.Cout(\timer[0]~26 ),
	.Q(timer[0]));
defparam \timer[0] .coord_x = 2;
defparam \timer[0] .coord_y = 12;
defparam \timer[0] .coord_z = 4;
defparam \timer[0] .mask = 16'h33CC;
defparam \timer[0] .modeMux = 1'b0;
defparam \timer[0] .FeedbackMux = 1'b0;
defparam \timer[0] .ShiftMux = 1'b0;
defparam \timer[0] .BypassEn = 1'b1;
defparam \timer[0] .CarryEnb = 1'b0;

alta_slice \timer[10] (
	.A(timer[10]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[9]~44 ),
	.Qin(timer[10]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y19_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y19_GND),
	.LutOut(\timer[10]~45_combout ),
	.Cout(\timer[10]~46 ),
	.Q(timer[10]));
defparam \timer[10] .coord_x = 2;
defparam \timer[10] .coord_y = 12;
defparam \timer[10] .coord_z = 14;
defparam \timer[10] .mask = 16'hA50A;
defparam \timer[10] .modeMux = 1'b1;
defparam \timer[10] .FeedbackMux = 1'b0;
defparam \timer[10] .ShiftMux = 1'b0;
defparam \timer[10] .BypassEn = 1'b1;
defparam \timer[10] .CarryEnb = 1'b0;

alta_slice \timer[11] (
	.A(timer[11]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[10]~46 ),
	.Qin(timer[11]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y19_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y19_GND),
	.LutOut(\timer[11]~47_combout ),
	.Cout(\timer[11]~48 ),
	.Q(timer[11]));
defparam \timer[11] .coord_x = 2;
defparam \timer[11] .coord_y = 12;
defparam \timer[11] .coord_z = 15;
defparam \timer[11] .mask = 16'h5A5F;
defparam \timer[11] .modeMux = 1'b1;
defparam \timer[11] .FeedbackMux = 1'b0;
defparam \timer[11] .ShiftMux = 1'b0;
defparam \timer[11] .BypassEn = 1'b1;
defparam \timer[11] .CarryEnb = 1'b0;

alta_slice \timer[12] (
	.A(timer[12]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[11]~48 ),
	.Qin(timer[12]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y18_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y18_GND),
	.LutOut(\timer[12]~49_combout ),
	.Cout(\timer[12]~50 ),
	.Q(timer[12]));
defparam \timer[12] .coord_x = 2;
defparam \timer[12] .coord_y = 11;
defparam \timer[12] .coord_z = 0;
defparam \timer[12] .mask = 16'hA50A;
defparam \timer[12] .modeMux = 1'b1;
defparam \timer[12] .FeedbackMux = 1'b0;
defparam \timer[12] .ShiftMux = 1'b0;
defparam \timer[12] .BypassEn = 1'b1;
defparam \timer[12] .CarryEnb = 1'b0;

alta_slice \timer[13] (
	.A(timer[13]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[12]~50 ),
	.Qin(timer[13]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y18_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y18_GND),
	.LutOut(\timer[13]~51_combout ),
	.Cout(\timer[13]~52 ),
	.Q(timer[13]));
defparam \timer[13] .coord_x = 2;
defparam \timer[13] .coord_y = 11;
defparam \timer[13] .coord_z = 1;
defparam \timer[13] .mask = 16'h5A5F;
defparam \timer[13] .modeMux = 1'b1;
defparam \timer[13] .FeedbackMux = 1'b0;
defparam \timer[13] .ShiftMux = 1'b0;
defparam \timer[13] .BypassEn = 1'b1;
defparam \timer[13] .CarryEnb = 1'b0;

alta_slice \timer[14] (
	.A(vcc),
	.B(timer[14]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[13]~52 ),
	.Qin(timer[14]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y18_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y18_GND),
	.LutOut(\timer[14]~53_combout ),
	.Cout(\timer[14]~54 ),
	.Q(timer[14]));
defparam \timer[14] .coord_x = 2;
defparam \timer[14] .coord_y = 11;
defparam \timer[14] .coord_z = 2;
defparam \timer[14] .mask = 16'hC30C;
defparam \timer[14] .modeMux = 1'b1;
defparam \timer[14] .FeedbackMux = 1'b0;
defparam \timer[14] .ShiftMux = 1'b0;
defparam \timer[14] .BypassEn = 1'b1;
defparam \timer[14] .CarryEnb = 1'b0;

alta_slice \timer[15] (
	.A(vcc),
	.B(timer[15]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[14]~54 ),
	.Qin(timer[15]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y18_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y18_GND),
	.LutOut(\timer[15]~55_combout ),
	.Cout(\timer[15]~56 ),
	.Q(timer[15]));
defparam \timer[15] .coord_x = 2;
defparam \timer[15] .coord_y = 11;
defparam \timer[15] .coord_z = 3;
defparam \timer[15] .mask = 16'h3C3F;
defparam \timer[15] .modeMux = 1'b1;
defparam \timer[15] .FeedbackMux = 1'b0;
defparam \timer[15] .ShiftMux = 1'b0;
defparam \timer[15] .BypassEn = 1'b1;
defparam \timer[15] .CarryEnb = 1'b0;

alta_slice \timer[16] (
	.A(vcc),
	.B(timer[16]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[15]~56 ),
	.Qin(timer[16]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y18_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y18_GND),
	.LutOut(\timer[16]~57_combout ),
	.Cout(\timer[16]~58 ),
	.Q(timer[16]));
defparam \timer[16] .coord_x = 2;
defparam \timer[16] .coord_y = 11;
defparam \timer[16] .coord_z = 4;
defparam \timer[16] .mask = 16'hC30C;
defparam \timer[16] .modeMux = 1'b1;
defparam \timer[16] .FeedbackMux = 1'b0;
defparam \timer[16] .ShiftMux = 1'b0;
defparam \timer[16] .BypassEn = 1'b1;
defparam \timer[16] .CarryEnb = 1'b0;

alta_slice \timer[17] (
	.A(timer[17]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[16]~58 ),
	.Qin(timer[17]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y18_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y18_GND),
	.LutOut(\timer[17]~59_combout ),
	.Cout(\timer[17]~60 ),
	.Q(timer[17]));
defparam \timer[17] .coord_x = 2;
defparam \timer[17] .coord_y = 11;
defparam \timer[17] .coord_z = 5;
defparam \timer[17] .mask = 16'h5A5F;
defparam \timer[17] .modeMux = 1'b1;
defparam \timer[17] .FeedbackMux = 1'b0;
defparam \timer[17] .ShiftMux = 1'b0;
defparam \timer[17] .BypassEn = 1'b1;
defparam \timer[17] .CarryEnb = 1'b0;

alta_slice \timer[18] (
	.A(vcc),
	.B(timer[18]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[17]~60 ),
	.Qin(timer[18]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y18_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y18_GND),
	.LutOut(\timer[18]~61_combout ),
	.Cout(\timer[18]~62 ),
	.Q(timer[18]));
defparam \timer[18] .coord_x = 2;
defparam \timer[18] .coord_y = 11;
defparam \timer[18] .coord_z = 6;
defparam \timer[18] .mask = 16'hC30C;
defparam \timer[18] .modeMux = 1'b1;
defparam \timer[18] .FeedbackMux = 1'b0;
defparam \timer[18] .ShiftMux = 1'b0;
defparam \timer[18] .BypassEn = 1'b1;
defparam \timer[18] .CarryEnb = 1'b0;

alta_slice \timer[19] (
	.A(timer[19]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[18]~62 ),
	.Qin(timer[19]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y18_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y18_GND),
	.LutOut(\timer[19]~63_combout ),
	.Cout(\timer[19]~64 ),
	.Q(timer[19]));
defparam \timer[19] .coord_x = 2;
defparam \timer[19] .coord_y = 11;
defparam \timer[19] .coord_z = 7;
defparam \timer[19] .mask = 16'h5A5F;
defparam \timer[19] .modeMux = 1'b1;
defparam \timer[19] .FeedbackMux = 1'b0;
defparam \timer[19] .ShiftMux = 1'b0;
defparam \timer[19] .BypassEn = 1'b1;
defparam \timer[19] .CarryEnb = 1'b0;

alta_slice \timer[1] (
	.A(timer[1]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[0]~26 ),
	.Qin(timer[1]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y19_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y19_GND),
	.LutOut(\timer[1]~27_combout ),
	.Cout(\timer[1]~28 ),
	.Q(timer[1]));
defparam \timer[1] .coord_x = 2;
defparam \timer[1] .coord_y = 12;
defparam \timer[1] .coord_z = 5;
defparam \timer[1] .mask = 16'h5A5F;
defparam \timer[1] .modeMux = 1'b1;
defparam \timer[1] .FeedbackMux = 1'b0;
defparam \timer[1] .ShiftMux = 1'b0;
defparam \timer[1] .BypassEn = 1'b1;
defparam \timer[1] .CarryEnb = 1'b0;

alta_slice \timer[20] (
	.A(vcc),
	.B(timer[20]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[19]~64 ),
	.Qin(timer[20]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y18_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y18_GND),
	.LutOut(\timer[20]~65_combout ),
	.Cout(\timer[20]~66 ),
	.Q(timer[20]));
defparam \timer[20] .coord_x = 2;
defparam \timer[20] .coord_y = 11;
defparam \timer[20] .coord_z = 8;
defparam \timer[20] .mask = 16'hC30C;
defparam \timer[20] .modeMux = 1'b1;
defparam \timer[20] .FeedbackMux = 1'b0;
defparam \timer[20] .ShiftMux = 1'b0;
defparam \timer[20] .BypassEn = 1'b1;
defparam \timer[20] .CarryEnb = 1'b0;

alta_slice \timer[21] (
	.A(vcc),
	.B(timer[21]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[20]~66 ),
	.Qin(timer[21]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y18_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y18_GND),
	.LutOut(\timer[21]~67_combout ),
	.Cout(\timer[21]~68 ),
	.Q(timer[21]));
defparam \timer[21] .coord_x = 2;
defparam \timer[21] .coord_y = 11;
defparam \timer[21] .coord_z = 9;
defparam \timer[21] .mask = 16'h3C3F;
defparam \timer[21] .modeMux = 1'b1;
defparam \timer[21] .FeedbackMux = 1'b0;
defparam \timer[21] .ShiftMux = 1'b0;
defparam \timer[21] .BypassEn = 1'b1;
defparam \timer[21] .CarryEnb = 1'b0;

alta_slice \timer[22] (
	.A(vcc),
	.B(timer[22]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[21]~68 ),
	.Qin(timer[22]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y18_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y18_GND),
	.LutOut(\timer[22]~69_combout ),
	.Cout(\timer[22]~70 ),
	.Q(timer[22]));
defparam \timer[22] .coord_x = 2;
defparam \timer[22] .coord_y = 11;
defparam \timer[22] .coord_z = 10;
defparam \timer[22] .mask = 16'hC30C;
defparam \timer[22] .modeMux = 1'b1;
defparam \timer[22] .FeedbackMux = 1'b0;
defparam \timer[22] .ShiftMux = 1'b0;
defparam \timer[22] .BypassEn = 1'b1;
defparam \timer[22] .CarryEnb = 1'b0;

alta_slice \timer[23] (
	.A(timer[23]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[22]~70 ),
	.Qin(timer[23]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y18_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y18_GND),
	.LutOut(\timer[23]~71_combout ),
	.Cout(\timer[23]~72 ),
	.Q(timer[23]));
defparam \timer[23] .coord_x = 2;
defparam \timer[23] .coord_y = 11;
defparam \timer[23] .coord_z = 11;
defparam \timer[23] .mask = 16'h5A5F;
defparam \timer[23] .modeMux = 1'b1;
defparam \timer[23] .FeedbackMux = 1'b0;
defparam \timer[23] .ShiftMux = 1'b0;
defparam \timer[23] .BypassEn = 1'b1;
defparam \timer[23] .CarryEnb = 1'b0;

alta_slice \timer[24] (
	.A(vcc),
	.B(timer[24]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[23]~72 ),
	.Qin(timer[24]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y18_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y18_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y18_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y18_GND),
	.LutOut(\timer[24]~73_combout ),
	.Cout(),
	.Q(timer[24]));
defparam \timer[24] .coord_x = 2;
defparam \timer[24] .coord_y = 11;
defparam \timer[24] .coord_z = 12;
defparam \timer[24] .mask = 16'hC3C3;
defparam \timer[24] .modeMux = 1'b1;
defparam \timer[24] .FeedbackMux = 1'b0;
defparam \timer[24] .ShiftMux = 1'b0;
defparam \timer[24] .BypassEn = 1'b1;
defparam \timer[24] .CarryEnb = 1'b1;

alta_slice \timer[2] (
	.A(vcc),
	.B(timer[2]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[1]~28 ),
	.Qin(timer[2]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y19_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y19_GND),
	.LutOut(\timer[2]~29_combout ),
	.Cout(\timer[2]~30 ),
	.Q(timer[2]));
defparam \timer[2] .coord_x = 2;
defparam \timer[2] .coord_y = 12;
defparam \timer[2] .coord_z = 6;
defparam \timer[2] .mask = 16'hC30C;
defparam \timer[2] .modeMux = 1'b1;
defparam \timer[2] .FeedbackMux = 1'b0;
defparam \timer[2] .ShiftMux = 1'b0;
defparam \timer[2] .BypassEn = 1'b1;
defparam \timer[2] .CarryEnb = 1'b0;

alta_slice \timer[3] (
	.A(timer[3]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[2]~30 ),
	.Qin(timer[3]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y19_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y19_GND),
	.LutOut(\timer[3]~31_combout ),
	.Cout(\timer[3]~32 ),
	.Q(timer[3]));
defparam \timer[3] .coord_x = 2;
defparam \timer[3] .coord_y = 12;
defparam \timer[3] .coord_z = 7;
defparam \timer[3] .mask = 16'h5A5F;
defparam \timer[3] .modeMux = 1'b1;
defparam \timer[3] .FeedbackMux = 1'b0;
defparam \timer[3] .ShiftMux = 1'b0;
defparam \timer[3] .BypassEn = 1'b1;
defparam \timer[3] .CarryEnb = 1'b0;

alta_slice \timer[4] (
	.A(vcc),
	.B(timer[4]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[3]~32 ),
	.Qin(timer[4]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y19_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y19_GND),
	.LutOut(\timer[4]~33_combout ),
	.Cout(\timer[4]~34 ),
	.Q(timer[4]));
defparam \timer[4] .coord_x = 2;
defparam \timer[4] .coord_y = 12;
defparam \timer[4] .coord_z = 8;
defparam \timer[4] .mask = 16'hC30C;
defparam \timer[4] .modeMux = 1'b1;
defparam \timer[4] .FeedbackMux = 1'b0;
defparam \timer[4] .ShiftMux = 1'b0;
defparam \timer[4] .BypassEn = 1'b1;
defparam \timer[4] .CarryEnb = 1'b0;

alta_slice \timer[5] (
	.A(vcc),
	.B(timer[5]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[4]~34 ),
	.Qin(timer[5]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y19_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y19_GND),
	.LutOut(\timer[5]~35_combout ),
	.Cout(\timer[5]~36 ),
	.Q(timer[5]));
defparam \timer[5] .coord_x = 2;
defparam \timer[5] .coord_y = 12;
defparam \timer[5] .coord_z = 9;
defparam \timer[5] .mask = 16'h3C3F;
defparam \timer[5] .modeMux = 1'b1;
defparam \timer[5] .FeedbackMux = 1'b0;
defparam \timer[5] .ShiftMux = 1'b0;
defparam \timer[5] .BypassEn = 1'b1;
defparam \timer[5] .CarryEnb = 1'b0;

alta_slice \timer[6] (
	.A(vcc),
	.B(timer[6]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[5]~36 ),
	.Qin(timer[6]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y19_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y19_GND),
	.LutOut(\timer[6]~37_combout ),
	.Cout(\timer[6]~38 ),
	.Q(timer[6]));
defparam \timer[6] .coord_x = 2;
defparam \timer[6] .coord_y = 12;
defparam \timer[6] .coord_z = 10;
defparam \timer[6] .mask = 16'hC30C;
defparam \timer[6] .modeMux = 1'b1;
defparam \timer[6] .FeedbackMux = 1'b0;
defparam \timer[6] .ShiftMux = 1'b0;
defparam \timer[6] .BypassEn = 1'b1;
defparam \timer[6] .CarryEnb = 1'b0;

alta_slice \timer[7] (
	.A(timer[7]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[6]~38 ),
	.Qin(timer[7]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y19_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y19_GND),
	.LutOut(\timer[7]~39_combout ),
	.Cout(\timer[7]~40 ),
	.Q(timer[7]));
defparam \timer[7] .coord_x = 2;
defparam \timer[7] .coord_y = 12;
defparam \timer[7] .coord_z = 11;
defparam \timer[7] .mask = 16'h5A5F;
defparam \timer[7] .modeMux = 1'b1;
defparam \timer[7] .FeedbackMux = 1'b0;
defparam \timer[7] .ShiftMux = 1'b0;
defparam \timer[7] .BypassEn = 1'b1;
defparam \timer[7] .CarryEnb = 1'b0;

alta_slice \timer[8] (
	.A(vcc),
	.B(timer[8]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[7]~40 ),
	.Qin(timer[8]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y19_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y19_GND),
	.LutOut(\timer[8]~41_combout ),
	.Cout(\timer[8]~42 ),
	.Q(timer[8]));
defparam \timer[8] .coord_x = 2;
defparam \timer[8] .coord_y = 12;
defparam \timer[8] .coord_z = 12;
defparam \timer[8] .mask = 16'hC30C;
defparam \timer[8] .modeMux = 1'b1;
defparam \timer[8] .FeedbackMux = 1'b0;
defparam \timer[8] .ShiftMux = 1'b0;
defparam \timer[8] .BypassEn = 1'b1;
defparam \timer[8] .CarryEnb = 1'b0;

alta_slice \timer[9] (
	.A(vcc),
	.B(timer[9]),
	.C(vcc),
	.D(vcc),
	.Cin(\timer[8]~42 ),
	.Qin(timer[9]),
	.Clk(\clk~inputclkctrl_outclk_X25_Y19_SIG_VCC ),
	.AsyncReset(AsyncReset_X25_Y19_GND),
	.SyncReset(\alt_pll_inst|altpll_component|auto_generated|locked~combout__SyncReset_X25_Y19_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X25_Y19_GND),
	.LutOut(\timer[9]~43_combout ),
	.Cout(\timer[9]~44 ),
	.Q(timer[9]));
defparam \timer[9] .coord_x = 2;
defparam \timer[9] .coord_y = 12;
defparam \timer[9] .coord_z = 13;
defparam \timer[9] .mask = 16'h3C3F;
defparam \timer[9] .modeMux = 1'b1;
defparam \timer[9] .FeedbackMux = 1'b0;
defparam \timer[9] .ShiftMux = 1'b0;
defparam \timer[9] .BypassEn = 1'b1;
defparam \timer[9] .CarryEnb = 1'b0;

alta_slice \~QIC_CREATED_GND~I (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\~QIC_CREATED_GND~I_combout ),
	.Cout(),
	.Q());
defparam \~QIC_CREATED_GND~I .coord_x = 6;
defparam \~QIC_CREATED_GND~I .coord_y = 10;
defparam \~QIC_CREATED_GND~I .coord_z = 12;
defparam \~QIC_CREATED_GND~I .mask = 16'h0000;
defparam \~QIC_CREATED_GND~I .modeMux = 1'b0;
defparam \~QIC_CREATED_GND~I .FeedbackMux = 1'b0;
defparam \~QIC_CREATED_GND~I .ShiftMux = 1'b0;
defparam \~QIC_CREATED_GND~I .BypassEn = 1'b0;
defparam \~QIC_CREATED_GND~I .CarryEnb = 1'b1;

endmodule
